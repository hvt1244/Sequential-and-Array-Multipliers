
module Add_half_0 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2047 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_0 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_0 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2047 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2046 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2045 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1023 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2046 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2045 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2044 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2043 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1022 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2044 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2043 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2042 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CND2X1 U2 ( .A(n1), .B(a), .Z(n4) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX2 U4 ( .A(b), .Z(n1) );
  CND2X1 U5 ( .A(b), .B(n2), .Z(n3) );
  CIVX2 U6 ( .A(a), .Z(n2) );
endmodule


module Add_half_2041 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1021 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2042 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2041 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_0 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n4, n1, n2;

  CANR2X2 U3 ( .A(c_out01), .B(c_in2), .C(n2), .D(c_out00), .Z(n4) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n4), .Z(c_out2) );
  Add_full_0 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0)
         );
  Add_full_1023 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1022 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1021 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n4), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n4), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_2040 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2039 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1020 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2040 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2039 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2038 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2037 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1019 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2038 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2037 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2036 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2035 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1018 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2036 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2035 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2034 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2033 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1017 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2034 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2033 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_255 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_1020 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1019 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1018 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1017 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_2032 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2031 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1016 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2032 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2031 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2030 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2029 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1015 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2030 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2029 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2028 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2027 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1014 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2028 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2027 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2026 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2025 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1013 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2026 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2025 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_254 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_1016 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1015 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1014 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1013 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_2024 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2023 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1012 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2024 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2023 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2022 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2021 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1011 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2022 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2021 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2020 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2019 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1010 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2020 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2019 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2018 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2017 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1009 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2018 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2017 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_253 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_1012 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1011 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1010 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1009 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_0 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n4, n1, n2, n3, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n5), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n5), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_0 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_255 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_254 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_253 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n5), .Z(n4) );
  CNIVXL U4 ( .A(n4), .Z(n3) );
  CAOR2XL U5 ( .A(s44[1]), .B(n2), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2XL U6 ( .A(s44[0]), .B(n2), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CIVX2 U7 ( .A(n4), .Z(n1) );
  CIVXL U11 ( .A(n3), .Z(n2) );
  CIVX2 U12 ( .A(c_in4), .Z(n5) );
endmodule


module Add_half_2016 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2015 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1008 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2016 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2015 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2014 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2013 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1007 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2014 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2013 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2012 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2011 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1006 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2012 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2011 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2010 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2009 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1005 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2010 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2009 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_252 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n5,
         n6;

  CAOR2X1 U6 ( .A(s4), .B(n3), .C(s3), .D(n6), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  Add_full_1008 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1007 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1006 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1005 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n5), .Z(n6) );
  COND2X1 U4 ( .A(n1), .B(n6), .C(n2), .D(n3), .Z(c_out2) );
  CIVX2 U5 ( .A(c_out10), .Z(n2) );
  CIVX2 U8 ( .A(c_out11), .Z(n1) );
  CIVX2 U9 ( .A(n6), .Z(n3) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_2008 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2007 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1004 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2008 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2007 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2006 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2005 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1003 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2006 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2005 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2004 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2003 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1002 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2004 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2003 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2002 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2001 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1001 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2002 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2001 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_251 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_1004 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1003 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1002 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1001 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_2000 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1999 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1000 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2000 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1999 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1998 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1997 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_999 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1998 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1997 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1996 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1995 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_998 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1996 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1995 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1994 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1993 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_997 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1994 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1993 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_250 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_1000 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_999 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_998 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_997 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1992 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1991 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_996 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1992 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1991 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1990 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1989 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_995 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1990 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1989 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1988 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1987 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_994 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1988 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1987 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1986 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1985 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_993 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1986 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1985 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_249 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_996 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_995 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_994 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_993 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_63 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_252 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_251 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_250 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_249 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1984 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1983 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_992 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1984 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1983 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1982 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1981 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_991 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1982 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1981 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1980 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1979 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_990 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1980 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1979 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1978 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1977 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_989 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1978 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1977 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_248 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_992 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_991 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_990 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_989 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1976 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1975 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_988 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1976 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1975 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1974 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1973 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_987 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1974 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1973 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1972 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1971 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_986 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1972 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1971 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1970 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1969 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_985 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1970 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1969 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_247 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_988 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_987 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_986 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_985 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1968 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1967 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_984 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1968 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1967 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1966 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1965 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_983 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1966 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1965 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1964 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1963 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_982 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1964 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1963 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1962 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1961 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_981 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1962 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1961 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_246 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_984 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_983 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_982 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_981 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1960 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1959 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_980 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1960 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1959 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1958 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1957 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_979 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1958 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1957 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1956 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1955 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_978 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1956 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1955 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1954 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1953 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_977 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1954 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1953 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_245 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_980 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_979 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_978 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_977 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_62 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_248 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_247 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_246 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_245 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1952 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1951 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_976 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1952 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1951 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1950 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1949 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_975 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1950 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1949 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1948 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1947 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_974 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1948 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1947 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1946 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1945 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_973 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1946 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1945 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_244 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_976 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_975 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_974 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_973 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1944 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1943 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_972 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1944 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1943 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1942 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1941 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_971 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1942 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1941 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1940 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1939 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_970 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1940 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1939 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1938 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1937 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_969 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1938 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1937 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_243 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_972 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_971 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_970 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_969 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1936 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1935 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_968 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1936 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1935 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1934 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1933 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_967 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1934 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1933 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1932 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1931 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_966 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1932 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1931 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1930 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1929 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_965 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1930 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1929 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_242 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_968 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_967 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_966 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_965 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1928 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1927 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_964 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1928 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1927 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1926 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1925 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_963 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1926 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1925 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1924 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1923 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_962 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1924 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1923 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1922 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1921 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_961 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1922 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1921 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_241 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_964 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_963 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_962 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_961 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U5 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_61 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_244 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_243 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_242 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_241 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2XL U5 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CIVX2 U6 ( .A(n3), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_0 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n4, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n3), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n3), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n3), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n3), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n2), .C(c_out810), .D(n1), .Z(c_out8) );
  bit4_0 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_63 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_62 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_61 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CANR2X1 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n3), .Z(n4) );
  CANR2X1 U4 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n3), .Z(n1) );
  CAOR2XL U5 ( .A(s84[3]), .B(n2), .C(s83[3]), .D(n1), .Z(sum8[7]) );
  CAOR2XL U6 ( .A(s84[0]), .B(n2), .C(s83[0]), .D(n1), .Z(sum8[4]) );
  CAOR2XL U7 ( .A(s84[1]), .B(n2), .C(s83[1]), .D(n1), .Z(sum8[5]) );
  CAOR2XL U8 ( .A(s84[2]), .B(n2), .C(s83[2]), .D(n1), .Z(sum8[6]) );
  CIVX2 U9 ( .A(n4), .Z(n2) );
  CIVX2 U15 ( .A(c_in8), .Z(n3) );
endmodule


module Add_half_1920 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1919 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CEOX1 U2 ( .A(b), .B(n1), .Z(sum) );
  CAN2X1 U3 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_960 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1920 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1919 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1918 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1917 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_959 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1918 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1917 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1916 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1915 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_958 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1916 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1915 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1914 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1913 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_957 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1914 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1913 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_240 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_960 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_959 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_958 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_957 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1912 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1911 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_956 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1912 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1911 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1910 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1909 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_955 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1910 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1909 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1908 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1907 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_954 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1908 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1907 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1906 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1905 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_953 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1906 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1905 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_239 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_956 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_955 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_954 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_953 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1904 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1903 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_952 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1904 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1903 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1902 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1901 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_951 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1902 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1901 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1900 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1899 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_950 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1900 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1899 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1898 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1897 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_949 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1898 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1897 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_238 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_952 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_951 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_950 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_949 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1896 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1895 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_948 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1896 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1895 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1894 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1893 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_947 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1894 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1893 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1892 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1891 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_946 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1892 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1891 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1890 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1889 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_945 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1890 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1889 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_237 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_948 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_947 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_946 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_945 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_60 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n3), .C(s43[1]), .D(n6), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n3), .C(s43[0]), .D(n6), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n5), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n5), .Z(sum4[0]) );
  bit2_240 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_239 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_238 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_237 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n5), .Z(n6) );
  COND2X1 U4 ( .A(n1), .B(n6), .C(n2), .D(n3), .Z(c_out4) );
  CIVX2 U5 ( .A(c_out410), .Z(n2) );
  CIVX2 U10 ( .A(c_out411), .Z(n1) );
  CIVX2 U11 ( .A(n6), .Z(n3) );
  CIVX2 U12 ( .A(c_in4), .Z(n5) );
endmodule


module Add_half_1888 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1887 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_944 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1888 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1887 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1886 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1885 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_943 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1886 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1885 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1884 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1883 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_942 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1884 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1883 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1882 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1881 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_941 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1882 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1881 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_236 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_944 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_943 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_942 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_941 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1880 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1879 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_940 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1880 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1879 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1878 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1877 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_939 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1878 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1877 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1876 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1875 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_938 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1876 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1875 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1874 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1873 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_937 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1874 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1873 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_235 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_940 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_939 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_938 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_937 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1872 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1871 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_936 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1872 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1871 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1870 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1869 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_935 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1870 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1869 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1868 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1867 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_934 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1868 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1867 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1866 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1865 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_933 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1866 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1865 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_234 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_936 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_935 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_934 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_933 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1864 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1863 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_932 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1864 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1863 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1862 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1861 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_931 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1862 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1861 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1860 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1859 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_930 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1860 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1859 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1858 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1857 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_929 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1858 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1857 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_233 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_932 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_931 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_930 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_929 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_59 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_236 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_235 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_234 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_233 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2XL U3 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2XL U4 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CANR2X2 U5 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(n3), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1856 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1855 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_928 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1856 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1855 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1854 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1853 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_927 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1854 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1853 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1852 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1851 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_926 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1852 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1851 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1850 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1849 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_925 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1850 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1849 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_232 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_928 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_927 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_926 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_925 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1848 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1847 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_924 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1848 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1847 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1846 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1845 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_923 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1846 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1845 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1844 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1843 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_922 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1844 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1843 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1842 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1841 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_921 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1842 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1841 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_231 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_924 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_923 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_922 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_921 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1840 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1839 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_920 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1840 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1839 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1838 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1837 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_919 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1838 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1837 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1836 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1835 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_918 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1836 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1835 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1834 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1833 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_917 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1834 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1833 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_230 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_920 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_919 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_918 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_917 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1832 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1831 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_916 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1832 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1831 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1830 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1829 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_915 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1830 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1829 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1828 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1827 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_914 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1828 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1827 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1826 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1825 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_913 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1826 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1825 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_229 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_916 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_915 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_914 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_913 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_58 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_232 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_231 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_230 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_229 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1824 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1823 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_912 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1824 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1823 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1822 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1821 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_911 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1822 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1821 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1820 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1819 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_910 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1820 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1819 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1818 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1817 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_909 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1818 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1817 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_228 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_912 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_911 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_910 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_909 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1816 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1815 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_908 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1816 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1815 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1814 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1813 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_907 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1814 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1813 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1812 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1811 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_906 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1812 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1811 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1810 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1809 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_905 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1810 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1809 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_227 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_908 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_907 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_906 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_905 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1808 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1807 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_904 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1808 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1807 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1806 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1805 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_903 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1806 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1805 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1804 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1803 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_902 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1804 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1803 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1802 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1801 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_901 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1802 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1801 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_226 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_904 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_903 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_902 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_901 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1800 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1799 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_900 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1800 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1799 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1798 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1797 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_899 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1798 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1797 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1796 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1795 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_898 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1796 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1795 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1794 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1793 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_897 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1794 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1793 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_225 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_900 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_899 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_898 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_897 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_57 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_228 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_227 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_226 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_225 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2XL U5 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CIVX2 U6 ( .A(n3), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_15 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n2), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n2), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n2), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n2), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n1), .C(c_out810), .D(n3), .Z(c_out8) );
  bit4_60 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_59 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_58 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_57 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVX2 U3 ( .A(n3), .Z(n1) );
  CANR2X2 U4 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n2), .Z(n3) );
  CAOR2XL U5 ( .A(s84[0]), .B(n1), .C(s83[0]), .D(n3), .Z(sum8[4]) );
  CAOR2XL U6 ( .A(s84[2]), .B(n1), .C(s83[2]), .D(n3), .Z(sum8[6]) );
  CAOR2XL U7 ( .A(s84[3]), .B(n1), .C(s83[3]), .D(n3), .Z(sum8[7]) );
  CAOR2XL U8 ( .A(s84[1]), .B(n1), .C(s83[1]), .D(n3), .Z(sum8[5]) );
  CIVX2 U9 ( .A(c_in8), .Z(n2) );
endmodule


module Add_half_1792 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVX1 U1 ( .A(a), .Z(n2) );
  CND2X1 U2 ( .A(b), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n1), .B(a), .Z(n4) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVX2 U5 ( .A(b), .Z(n1) );
  CAN2X1 U6 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1791 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_896 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1792 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1791 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1790 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1789 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_895 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1790 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1789 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1788 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1787 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_894 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1788 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1787 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1786 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1785 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_893 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1786 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1785 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_224 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_896 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_895 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_894 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_893 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1784 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1783 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_892 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1784 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1783 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1782 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1781 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_891 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1782 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1781 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1780 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1779 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_890 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1780 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1779 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1778 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1777 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_889 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1778 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1777 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_223 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_892 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_891 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_890 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_889 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1776 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1775 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_888 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1776 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1775 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1774 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1773 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_887 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1774 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1773 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1772 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1771 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_886 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1772 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1771 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1770 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1769 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_885 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1770 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1769 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_222 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_888 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_887 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_886 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_885 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1768 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1767 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_884 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1768 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1767 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1766 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1765 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_883 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1766 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1765 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1764 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1763 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_882 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1764 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1763 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1762 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1761 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_881 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1762 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1761 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_221 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_884 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_883 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_882 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_881 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_56 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_224 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_223 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_222 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_221 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1760 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1759 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_880 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1760 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1759 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1758 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1757 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_879 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1758 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1757 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1756 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1755 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_878 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1756 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1755 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1754 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1753 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_877 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1754 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1753 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_220 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_880 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_879 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_878 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_877 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1752 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1751 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_876 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1752 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1751 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1750 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1749 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_875 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1750 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1749 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1748 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1747 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_874 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1748 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1747 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1746 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1745 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_873 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1746 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1745 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_219 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_876 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_875 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_874 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_873 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1744 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1743 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_872 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1744 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1743 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1742 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1741 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_871 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1742 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1741 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1740 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1739 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_870 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1740 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1739 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1738 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1737 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_869 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1738 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1737 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_218 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  Add_full_872 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_871 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_870 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_869 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U8 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1736 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1735 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_868 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1736 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1735 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1734 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1733 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_867 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1734 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1733 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1732 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1731 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_866 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1732 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1731 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1730 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1729 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_865 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1730 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1729 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_217 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_868 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_867 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_866 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_865 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_55 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_220 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_219 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_218 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_217 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1728 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1727 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_864 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1728 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1727 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1726 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1725 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_863 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1726 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1725 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1724 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1723 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_862 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1724 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1723 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1722 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1721 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_861 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1722 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1721 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_216 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_864 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_863 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_862 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_861 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1720 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1719 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_860 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1720 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1719 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1718 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1717 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_859 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1718 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1717 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1716 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1715 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_858 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1716 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1715 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1714 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1713 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_857 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1714 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1713 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_215 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_860 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_859 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_858 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_857 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1712 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1711 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_856 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1712 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1711 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1710 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1709 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_855 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1710 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1709 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1708 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1707 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_854 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1708 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1707 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1706 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1705 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_853 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1706 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1705 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_214 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_856 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_855 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_854 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_853 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1704 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1703 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_852 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1704 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1703 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1702 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1701 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_851 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1702 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1701 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1700 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1699 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_850 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1700 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1699 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1698 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1697 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_849 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1698 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1697 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_213 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_852 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_851 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_850 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_849 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_54 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_216 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_215 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_214 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_213 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1696 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1695 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_848 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1696 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1695 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1694 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1693 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_847 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1694 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1693 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1692 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1691 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_846 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1692 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1691 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1690 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1689 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_845 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1690 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1689 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_212 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_848 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_847 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_846 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_845 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1688 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1687 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_844 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1688 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1687 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1686 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1685 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_843 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1686 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1685 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1684 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1683 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_842 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1684 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1683 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1682 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1681 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_841 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1682 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1681 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_211 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_844 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_843 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_842 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_841 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1680 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1679 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_840 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1680 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1679 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1678 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1677 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_839 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1678 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1677 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1676 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1675 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_838 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1676 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1675 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1674 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1673 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_837 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1674 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1673 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_210 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_840 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_839 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_838 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_837 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1672 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1671 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_836 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1672 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1671 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1670 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1669 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_835 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1670 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1669 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1668 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1667 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_834 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1668 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1667 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1666 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1665 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_833 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1666 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1665 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_209 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_836 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_835 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_834 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_833 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_53 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_212 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_211 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_210 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_209 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_14 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U6 ( .A(s84[3]), .B(n2), .C(s83[3]), .D(n1), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n2), .C(s83[2]), .D(n1), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n2), .C(s83[1]), .D(n1), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n2), .C(s83[0]), .D(n1), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n3), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n3), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n3), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n3), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n2), .C(c_out810), .D(n1), .Z(c_out8) );
  bit4_56 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_55 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_54 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_53 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CANR2X1 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n3), .Z(n5) );
  CNIVX1 U4 ( .A(n5), .Z(n1) );
  CIVX2 U5 ( .A(n5), .Z(n2) );
  CIVX2 U15 ( .A(c_in8), .Z(n3) );
endmodule


module Add_half_1664 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1663 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_832 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1664 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1663 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1662 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1661 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_831 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1662 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1661 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1660 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1659 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_830 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1660 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1659 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1658 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1657 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_829 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1658 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1657 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_208 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n2), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n2), .Z(c_out2) );
  Add_full_832 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_831 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_830 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_829 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n3), .Z(n1) );
  CANR2XL U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n3), .Z(n2) );
  CIVX2 U5 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_1656 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1655 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_828 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1656 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1655 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1654 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1653 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_827 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1654 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1653 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1652 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1651 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_826 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1652 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1651 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1650 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1649 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_825 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1650 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1649 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_207 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_828 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_827 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_826 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_825 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1648 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1647 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_824 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1648 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1647 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1646 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1645 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_823 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1646 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1645 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1644 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1643 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_822 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1644 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1643 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1642 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1641 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_821 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1642 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1641 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_206 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_824 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_823 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_822 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_821 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1640 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1639 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_820 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1640 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1639 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1638 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1637 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_819 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1638 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1637 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1636 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1635 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_818 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1636 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1635 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1634 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1633 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_817 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1634 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1633 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_205 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_820 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_819 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_818 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_817 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_52 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_208 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_207 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_206 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_205 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1632 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1631 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_816 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1632 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1631 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1630 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1629 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_815 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1630 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1629 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1628 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1627 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_814 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1628 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1627 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1626 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1625 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_813 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1626 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1625 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_204 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n5,
         n6;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n3), .C(c_out10), .D(n6), .Z(c_out2) );
  Add_full_816 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_815 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_814 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_813 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAN2X1 U3 ( .A(n1), .B(n2), .Z(n6) );
  CND2X1 U4 ( .A(c_out00), .B(n5), .Z(n2) );
  CND2X1 U5 ( .A(c_out01), .B(c_in2), .Z(n1) );
  CAOR2XL U6 ( .A(s4), .B(n3), .C(s3), .D(n6), .Z(sum2[1]) );
  CIVX2 U9 ( .A(n6), .Z(n3) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_1624 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1623 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_812 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1624 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1623 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1622 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1621 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_811 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1622 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1621 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1620 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1619 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_810 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1620 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1619 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1618 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1617 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_809 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1618 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1617 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_203 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_812 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_811 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_810 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_809 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1616 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1615 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_808 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1616 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1615 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1614 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1613 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_807 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1614 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1613 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1612 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1611 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_806 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1612 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1611 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1610 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1609 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_805 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1610 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1609 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_202 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_808 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_807 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_806 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_805 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1608 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1607 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_804 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1608 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1607 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1606 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1605 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_803 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1606 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1605 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1604 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1603 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_802 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1604 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1603 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1602 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1601 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_801 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1602 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1601 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_201 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_804 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_803 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_802 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_801 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_51 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_204 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_203 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_202 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_201 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1600 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1599 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_800 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1600 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1599 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1598 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1597 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_799 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1598 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1597 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1596 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1595 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_798 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1596 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1595 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1594 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1593 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_797 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1594 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1593 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_200 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_800 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_799 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_798 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_797 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1592 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1591 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_796 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1592 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1591 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1590 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1589 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_795 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1590 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1589 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1588 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1587 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_794 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1588 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1587 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1586 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1585 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_793 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1586 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1585 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_199 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_796 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_795 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_794 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_793 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1584 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1583 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_792 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1584 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1583 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1582 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1581 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_791 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1582 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1581 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1580 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1579 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_790 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1580 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1579 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1578 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1577 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_789 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1578 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1577 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_198 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_792 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_791 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_790 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_789 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1576 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1575 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_788 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1576 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1575 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1574 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1573 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_787 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1574 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1573 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1572 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1571 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_786 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1572 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1571 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1570 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1569 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_785 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1570 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1569 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_197 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_788 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_787 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_786 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_785 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_50 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_200 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_199 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_198 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_197 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1568 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1567 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_784 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1568 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1567 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1566 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1565 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_783 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1566 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1565 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1564 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1563 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_782 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1564 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1563 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1562 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1561 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_781 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1562 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1561 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_196 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_784 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_783 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_782 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_781 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1560 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1559 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_780 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1560 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1559 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1558 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1557 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_779 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1558 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1557 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1556 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1555 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_778 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1556 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1555 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1554 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1553 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_777 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1554 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1553 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_195 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_780 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_779 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_778 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_777 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1552 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1551 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_776 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1552 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1551 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1550 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1549 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_775 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1550 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1549 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1548 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1547 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_774 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1548 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1547 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1546 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1545 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_773 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1546 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1545 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_194 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_776 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_775 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_774 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_773 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1544 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1543 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_772 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1544 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1543 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1542 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1541 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_771 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1542 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1541 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1540 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1539 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_770 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1540 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1539 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1538 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1537 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_769 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1538 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1537 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_193 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_772 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_771 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_770 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_769 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_49 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_196 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_195 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_194 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_193 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2XL U5 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CIVX2 U6 ( .A(n3), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_13 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n3), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n3), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n3), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n3), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n1), .C(c_out810), .D(n2), .Z(c_out8) );
  bit4_52 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_51 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_50 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_49 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CAOR2X2 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n3), .Z(n1) );
  CIVX1 U4 ( .A(n1), .Z(n2) );
  CAOR2XL U5 ( .A(s84[0]), .B(n1), .C(s83[0]), .D(n2), .Z(sum8[4]) );
  CAOR2XL U6 ( .A(s84[1]), .B(n1), .C(s83[1]), .D(n2), .Z(sum8[5]) );
  CAOR2XL U7 ( .A(s84[2]), .B(n1), .C(s83[2]), .D(n2), .Z(sum8[6]) );
  CAOR2XL U8 ( .A(s84[3]), .B(n1), .C(s83[3]), .D(n2), .Z(sum8[7]) );
  CIVX2 U9 ( .A(c_in8), .Z(n3) );
endmodule


module bit16_0 ( sum16, c_out16, a16, b16, c_in16 );
  output [15:0] sum16;
  input [15:0] a16;
  input [15:0] b16;
  input c_in16;
  output c_out16;
  wire   c_out1600, c_out1601, c_out1610, c_out1611, n4, n1, n2, n3, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37;
  wire   [7:0] s161;
  wire   [7:0] s162;
  wire   [7:0] s163;
  wire   [7:0] s164;

  CAOR2X1 U8 ( .A(s162[7]), .B(c_in16), .C(s161[7]), .D(n37), .Z(sum16[7]) );
  CAOR2X1 U9 ( .A(s162[6]), .B(c_in16), .C(s161[6]), .D(n37), .Z(sum16[6]) );
  CAOR2X1 U10 ( .A(s162[5]), .B(c_in16), .C(s161[5]), .D(n37), .Z(sum16[5]) );
  CAOR2X1 U11 ( .A(s162[4]), .B(c_in16), .C(s161[4]), .D(n37), .Z(sum16[4]) );
  CAOR2X1 U12 ( .A(s162[3]), .B(c_in16), .C(s161[3]), .D(n37), .Z(sum16[3]) );
  CAOR2X1 U13 ( .A(s162[2]), .B(c_in16), .C(s161[2]), .D(n37), .Z(sum16[2]) );
  CAOR2X1 U14 ( .A(s162[1]), .B(c_in16), .C(s161[1]), .D(n37), .Z(sum16[1]) );
  CAOR2X1 U21 ( .A(s162[0]), .B(c_in16), .C(s161[0]), .D(n37), .Z(sum16[0]) );
  CAOR2X1 U22 ( .A(c_out1611), .B(n36), .C(c_out1610), .D(n5), .Z(c_out16) );
  bit8_0 A161 ( .sum8(s161), .c_out8(c_out1600), .a8({n28, n27, n26, n25, n24, 
        n23, n22, n21}), .b8({n8, n15, n14, n13, n12, n11, n10, n9}), .c_in8(
        1'b0) );
  bit8_15 A162 ( .sum8(s162), .c_out8(c_out1601), .a8({n28, n27, n26, n25, n24, 
        n23, n22, n21}), .b8({n8, n15, n14, n13, n12, n11, n10, n9}), .c_in8(
        1'b1) );
  bit8_14 A163 ( .sum8(s163), .c_out8(c_out1610), .a8({n35, n34, n33, n32, n31, 
        n30, n29, n6}), .b8({n20, n19, b16[13], n18, n7, n1, n17, n16}), 
        .c_in8(1'b0) );
  bit8_13 A164 ( .sum8(s164), .c_out8(c_out1611), .a8({n35, n34, n33, n32, n31, 
        n30, n29, n6}), .b8({n20, n19, b16[13], n18, n7, n1, n17, n16}), 
        .c_in8(1'b1) );
  CNIVX4 U3 ( .A(a16[8]), .Z(n6) );
  CNIVX2 U4 ( .A(a16[2]), .Z(n23) );
  CNIVX2 U5 ( .A(a16[4]), .Z(n25) );
  CNIVX2 U6 ( .A(b16[3]), .Z(n12) );
  CNIVX2 U7 ( .A(b16[6]), .Z(n15) );
  CNIVX1 U15 ( .A(b16[7]), .Z(n8) );
  CNIVX1 U16 ( .A(b16[11]), .Z(n7) );
  CNIVX2 U17 ( .A(b16[1]), .Z(n10) );
  CNIVX2 U18 ( .A(a16[1]), .Z(n22) );
  CNIVX2 U19 ( .A(b16[10]), .Z(n1) );
  CNIVXL U20 ( .A(n5), .Z(n2) );
  CNIVX4 U23 ( .A(b16[0]), .Z(n9) );
  CIVX2 U24 ( .A(n4), .Z(n36) );
  CANR2X1 U25 ( .A(c_out1601), .B(c_in16), .C(c_out1600), .D(n37), .Z(n4) );
  CNIVX2 U26 ( .A(b16[2]), .Z(n11) );
  CNIVX2 U27 ( .A(b16[4]), .Z(n13) );
  CANR2XL U28 ( .A(c_out1601), .B(c_in16), .C(c_out1600), .D(n37), .Z(n3) );
  CANR2XL U29 ( .A(c_out1601), .B(c_in16), .C(c_out1600), .D(n37), .Z(n5) );
  CNIVX3 U30 ( .A(b16[8]), .Z(n16) );
  CNIVX1 U31 ( .A(b16[5]), .Z(n14) );
  CNIVX2 U32 ( .A(b16[9]), .Z(n17) );
  CNIVX2 U33 ( .A(b16[12]), .Z(n18) );
  CNIVX2 U34 ( .A(a16[9]), .Z(n29) );
  CNIVX2 U35 ( .A(a16[5]), .Z(n26) );
  CNIVX2 U36 ( .A(a16[10]), .Z(n30) );
  CNIVX2 U37 ( .A(a16[6]), .Z(n27) );
  CNIVX2 U38 ( .A(a16[12]), .Z(n32) );
  CNIVX2 U39 ( .A(a16[3]), .Z(n24) );
  CNIVX1 U40 ( .A(b16[15]), .Z(n20) );
  CNIVX1 U41 ( .A(b16[14]), .Z(n19) );
  CNIVX4 U42 ( .A(a16[0]), .Z(n21) );
  CNIVX1 U43 ( .A(a16[15]), .Z(n35) );
  CNIVX1 U44 ( .A(a16[7]), .Z(n28) );
  CNIVX1 U45 ( .A(a16[11]), .Z(n31) );
  CNIVX1 U46 ( .A(a16[13]), .Z(n33) );
  CNIVX1 U47 ( .A(a16[14]), .Z(n34) );
  CAOR2XL U48 ( .A(s164[1]), .B(n36), .C(s163[1]), .D(n2), .Z(sum16[9]) );
  CAOR2XL U49 ( .A(s164[5]), .B(n36), .C(s163[5]), .D(n2), .Z(sum16[13]) );
  CAOR2XL U50 ( .A(s164[4]), .B(n36), .C(s163[4]), .D(n2), .Z(sum16[12]) );
  CAOR2XL U51 ( .A(s164[3]), .B(n36), .C(s163[3]), .D(n2), .Z(sum16[11]) );
  CAOR2XL U52 ( .A(s164[2]), .B(n36), .C(s163[2]), .D(n3), .Z(sum16[10]) );
  CAOR2XL U53 ( .A(s164[0]), .B(n36), .C(s163[0]), .D(n2), .Z(sum16[8]) );
  CAOR2XL U54 ( .A(s164[7]), .B(n36), .C(s163[7]), .D(n2), .Z(sum16[15]) );
  CAOR2XL U55 ( .A(s164[6]), .B(n36), .C(s163[6]), .D(n2), .Z(sum16[14]) );
  CIVX2 U56 ( .A(c_in16), .Z(n37) );
endmodule


module Add_half_1536 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1535 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_768 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1536 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1535 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1534 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1533 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_767 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1534 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1533 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1532 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1531 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_766 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1532 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1531 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1530 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVXL U1 ( .A(a), .Z(n1) );
  CENX1 U2 ( .A(b), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1529 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_765 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1530 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1529 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_192 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n5,
         n6;

  CAOR2X1 U6 ( .A(s4), .B(n3), .C(s3), .D(n6), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  Add_full_768 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_767 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_766 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_765 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n5), .Z(n6) );
  COND2X1 U4 ( .A(n1), .B(n6), .C(n2), .D(n3), .Z(c_out2) );
  CIVX2 U5 ( .A(c_out10), .Z(n2) );
  CIVX2 U8 ( .A(c_out11), .Z(n1) );
  CIVX2 U9 ( .A(n6), .Z(n3) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_1528 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1527 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_764 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1528 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1527 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1526 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1525 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_763 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1526 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1525 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1524 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1523 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_762 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1524 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1523 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1522 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1521 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_761 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1522 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1521 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_191 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_764 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_763 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_762 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_761 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X2 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1520 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1519 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_760 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1520 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1519 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1518 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1517 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_759 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1518 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1517 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1516 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1515 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_758 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1516 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1515 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1514 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1513 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_757 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1514 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1513 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_190 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_760 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_759 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_758 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_757 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1512 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1511 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_756 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1512 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1511 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1510 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1509 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_755 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1510 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1509 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1508 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1507 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_754 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1508 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1507 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1506 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1505 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_753 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1506 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1505 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_189 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_756 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_755 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_754 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_753 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_48 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_192 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_191 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_190 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_189 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2XL U5 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CIVX2 U6 ( .A(n3), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1504 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(b), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n1), .B(a), .Z(n4) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(b), .Z(n1) );
  CIVXL U5 ( .A(a), .Z(n2) );
  CAN2X1 U6 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1503 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_752 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1504 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1503 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1502 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1501 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_751 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1502 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1501 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1500 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1499 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_750 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1500 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1499 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1498 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1497 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_749 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1498 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1497 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_188 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n5,
         n6;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n3), .C(c_out10), .D(n6), .Z(c_out2) );
  Add_full_752 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_751 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_750 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_749 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAN2X1 U3 ( .A(n1), .B(n2), .Z(n6) );
  CND2X1 U4 ( .A(c_out01), .B(c_in2), .Z(n1) );
  CND2X1 U5 ( .A(c_out00), .B(n5), .Z(n2) );
  CAOR2XL U6 ( .A(s4), .B(n3), .C(s3), .D(n6), .Z(sum2[1]) );
  CIVX2 U9 ( .A(n6), .Z(n3) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_1496 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1495 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_748 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1496 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1495 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1494 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1493 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_747 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1494 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1493 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1492 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1491 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_746 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1492 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1491 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1490 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1489 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_745 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1490 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1489 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_187 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_748 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_747 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_746 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_745 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1488 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1487 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_744 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1488 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1487 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1486 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1485 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_743 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1486 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1485 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1484 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1483 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_742 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1484 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1483 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1482 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1481 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_741 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1482 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1481 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_186 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_744 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_743 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_742 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_741 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1480 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1479 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_740 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1480 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1479 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1478 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1477 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_739 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1478 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1477 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1476 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1475 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_738 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1476 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1475 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1474 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1473 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_737 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1474 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1473 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_185 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_740 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_739 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_738 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_737 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_47 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_188 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_187 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_186 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_185 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2XL U5 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CIVX2 U6 ( .A(n3), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1472 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX1 U1 ( .A(b), .B(n1), .Z(sum) );
  CIVX1 U2 ( .A(a), .Z(n1) );
  CAN2XL U3 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1471 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_736 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1472 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1471 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1470 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1469 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_735 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1470 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1469 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1468 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1467 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_734 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1468 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1467 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1466 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1465 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_733 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1466 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1465 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_184 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_736 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_735 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_734 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_733 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1464 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1463 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_732 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1464 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1463 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1462 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1461 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_731 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1462 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1461 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1460 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1459 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_730 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1460 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1459 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1458 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1457 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_729 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1458 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1457 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_183 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_732 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_731 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_730 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_729 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1456 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1455 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_728 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1456 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1455 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1454 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1453 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_727 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1454 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1453 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1452 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1451 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_726 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1452 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1451 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1450 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1449 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_725 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1450 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1449 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_182 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_728 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_727 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_726 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_725 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1448 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1447 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_724 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1448 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1447 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1446 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1445 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_723 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1446 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1445 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1444 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1443 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_722 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1444 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1443 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1442 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1441 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_721 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1442 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1441 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_181 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_724 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_723 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_722 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_721 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_46 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_184 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_183 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_182 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_181 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1440 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1439 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_720 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1440 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1439 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1438 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1437 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_719 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1438 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1437 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1436 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1435 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_718 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1436 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1435 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1434 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1433 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_717 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1434 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1433 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_180 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n2), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n2), .Z(c_out2) );
  Add_full_720 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_719 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_718 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_717 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n3), .Z(n2) );
  CIVX2 U5 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_1432 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1431 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_716 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1432 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1431 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1430 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1429 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_715 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1430 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1429 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1428 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1427 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_714 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1428 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1427 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1426 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1425 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_713 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1426 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1425 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_179 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_716 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_715 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_714 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_713 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1424 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1423 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_712 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1424 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1423 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1422 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1421 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_711 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1422 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1421 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1420 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1419 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_710 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1420 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1419 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1418 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1417 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_709 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1418 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1417 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_178 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_712 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_711 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_710 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_709 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1416 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1415 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_708 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1416 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1415 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1414 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1413 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_707 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1414 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1413 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1412 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1411 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_706 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1412 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1411 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1410 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1409 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_705 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1410 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1409 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_177 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_708 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_707 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_706 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_705 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_45 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_180 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_179 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_178 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_177 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2XL U5 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CIVX2 U6 ( .A(n3), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_12 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n5, n6;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n5), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n5), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n5), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n5), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n3), .C(c_out810), .D(n2), .Z(c_out8) );
  bit4_48 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_47 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_46 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_45 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CANR2X2 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n5), .Z(n6) );
  CAOR2XL U4 ( .A(s84[0]), .B(n3), .C(s83[0]), .D(n2), .Z(sum8[4]) );
  CAOR2XL U5 ( .A(s84[1]), .B(n3), .C(s83[1]), .D(n2), .Z(sum8[5]) );
  CAOR2XL U6 ( .A(s84[2]), .B(n3), .C(s83[2]), .D(n2), .Z(sum8[6]) );
  CAOR2XL U7 ( .A(s84[3]), .B(n3), .C(s83[3]), .D(n2), .Z(sum8[7]) );
  CIVXL U8 ( .A(n6), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n2) );
  CIVX2 U15 ( .A(n6), .Z(n3) );
  CIVX2 U16 ( .A(c_in8), .Z(n5) );
endmodule


module Add_half_1408 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1407 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_704 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1408 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1407 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1406 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1405 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_703 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1406 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1405 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1404 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1403 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_702 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1404 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1403 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1402 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1401 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_701 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1402 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1401 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_176 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_704 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_703 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_702 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_701 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X2 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1400 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1399 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_700 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1400 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1399 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1398 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1397 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_699 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1398 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1397 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1396 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1395 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_698 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1396 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1395 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1394 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1393 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_697 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1394 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1393 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_175 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_700 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_699 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_698 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_697 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1392 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1391 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_696 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1392 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1391 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1390 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1389 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_695 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1390 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1389 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1388 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1387 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_694 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1388 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1387 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1386 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1385 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_693 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1386 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1385 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_174 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_696 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_695 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_694 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_693 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1384 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1383 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_692 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1384 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1383 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1382 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1381 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_691 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1382 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1381 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1380 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1379 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_690 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1380 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1379 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1378 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1377 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_689 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1378 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1377 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_173 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_692 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_691 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_690 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_689 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_44 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n3), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n3), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n2), .Z(c_out4) );
  bit2_176 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_175 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_174 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_173 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n3), .Z(n5) );
  CIVDX1 U4 ( .A(n5), .Z0(n1), .Z1(n2) );
  CAOR2XL U5 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n2), .Z(sum4[3]) );
  CAOR2XL U6 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n2), .Z(sum4[2]) );
  CIVX2 U7 ( .A(c_in4), .Z(n3) );
endmodule


module Add_half_1376 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1375 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_688 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1376 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1375 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1374 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1373 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_687 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1374 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1373 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1372 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1371 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_686 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1372 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1371 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1370 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1369 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_685 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1370 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1369 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_172 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_688 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_687 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_686 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_685 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1368 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1367 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_684 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1368 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1367 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1366 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1365 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_683 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1366 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1365 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1364 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1363 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_682 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1364 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1363 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1362 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1361 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_681 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1362 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1361 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_171 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_684 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_683 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_682 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_681 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1360 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1359 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_680 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1360 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1359 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1358 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1357 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_679 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1358 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1357 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1356 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1355 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_678 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1356 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1355 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1354 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1353 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_677 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1354 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1353 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_170 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_680 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_679 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_678 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_677 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1352 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1351 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_676 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1352 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1351 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1350 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1349 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_675 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1350 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1349 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1348 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1347 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_674 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1348 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1347 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1346 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1345 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_673 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1346 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1345 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_169 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_676 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_675 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_674 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_673 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CAOR2XL U5 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_43 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_172 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_171 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_170 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_169 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1344 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1343 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_672 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1344 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1343 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1342 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1341 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_671 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1342 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1341 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1340 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1339 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_670 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1340 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1339 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1338 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1337 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_669 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1338 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1337 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_168 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_672 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_671 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_670 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_669 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1336 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1335 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_668 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1336 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1335 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1334 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1333 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_667 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1334 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1333 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1332 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1331 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_666 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1332 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1331 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1330 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1329 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_665 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1330 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1329 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_167 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_668 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_667 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_666 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_665 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1328 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1327 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_664 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1328 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1327 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1326 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1325 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_663 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1326 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1325 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1324 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1323 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_662 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1324 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1323 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1322 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1321 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_661 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1322 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1321 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_166 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_664 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_663 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_662 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_661 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1320 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1319 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_660 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1320 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1319 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1318 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1317 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_659 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1318 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1317 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1316 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1315 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_658 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1316 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1315 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1314 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1313 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_657 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1314 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1313 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_165 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_660 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_659 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_658 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_657 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_42 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_168 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_167 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_166 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_165 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2XL U5 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CIVX2 U6 ( .A(n3), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1312 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(b), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n1), .B(a), .Z(n4) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(b), .Z(n1) );
  CIVXL U5 ( .A(a), .Z(n2) );
  CAN2XL U6 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1311 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_656 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1312 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1311 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1310 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1309 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_655 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1310 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1309 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1308 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1307 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_654 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1308 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1307 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1306 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1305 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_653 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1306 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1305 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_164 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_656 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_655 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_654 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_653 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1304 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1303 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_652 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1304 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1303 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1302 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1301 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_651 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1302 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1301 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1300 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1299 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_650 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1300 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1299 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1298 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1297 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_649 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1298 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1297 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_163 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_652 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_651 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_650 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_649 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CAOR2XL U5 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1296 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1295 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_648 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1296 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1295 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1294 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1293 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_647 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1294 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1293 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1292 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1291 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_646 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1292 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1291 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1290 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1289 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_645 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1290 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1289 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_162 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_648 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_647 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_646 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_645 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1288 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1287 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_644 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1288 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1287 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1286 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1285 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_643 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1286 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1285 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1284 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1283 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_642 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1284 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1283 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1282 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1281 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_641 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1282 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1281 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_161 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_644 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_643 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_642 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_641 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_41 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n2), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n2), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n3), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n3), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n2), .Z(c_out4) );
  bit2_164 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_163 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_162 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_161 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVDX1 U3 ( .A(n5), .Z0(n1), .Z1(n2) );
  CANR2X1 U4 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n3), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n3) );
endmodule


module bit8_11 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n2), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n2), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n2), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n2), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n1), .C(c_out810), .D(n3), .Z(c_out8) );
  bit4_44 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_43 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_42 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_41 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CAOR2XL U3 ( .A(s84[3]), .B(n1), .C(s83[3]), .D(n3), .Z(sum8[7]) );
  CAOR2XL U4 ( .A(s84[2]), .B(n1), .C(s83[2]), .D(n3), .Z(sum8[6]) );
  CAOR2XL U5 ( .A(s84[1]), .B(n1), .C(s83[1]), .D(n3), .Z(sum8[5]) );
  CAOR2XL U6 ( .A(s84[0]), .B(n1), .C(s83[0]), .D(n3), .Z(sum8[4]) );
  CIVX2 U7 ( .A(n3), .Z(n1) );
  CANR2X2 U8 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n2), .Z(n3) );
  CIVX2 U9 ( .A(c_in8), .Z(n2) );
endmodule


module Add_half_1280 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVXL U1 ( .A(a), .Z(n1) );
  CENX1 U2 ( .A(b), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1279 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_640 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1280 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1279 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1278 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1277 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_639 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1278 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1277 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1276 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1275 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_638 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1276 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1275 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1274 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1273 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_637 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1274 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1273 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_160 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_640 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_639 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_638 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_637 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1272 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1271 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_636 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1272 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1271 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1270 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1269 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_635 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1270 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1269 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1268 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1267 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_634 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1268 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1267 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1266 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1265 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_633 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1266 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1265 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_159 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_636 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_635 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_634 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_633 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1264 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1263 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_632 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1264 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1263 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1262 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1261 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_631 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1262 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1261 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1260 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1259 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_630 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1260 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1259 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1258 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1257 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_629 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1258 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1257 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_158 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_632 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_631 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_630 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_629 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1256 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1255 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_628 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1256 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1255 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1254 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1253 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_627 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1254 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1253 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1252 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1251 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_626 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1252 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1251 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1250 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1249 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_625 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1250 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1249 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_157 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_628 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_627 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_626 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_625 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_40 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_160 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_159 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_158 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_157 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1248 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1247 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_624 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1248 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1247 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1246 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1245 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_623 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1246 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1245 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1244 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1243 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_622 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1244 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1243 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1242 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1241 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_621 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1242 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1241 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_156 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_624 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_623 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_622 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_621 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1240 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1239 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_620 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1240 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1239 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1238 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1237 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_619 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1238 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1237 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1236 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1235 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_618 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1236 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1235 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1234 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1233 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_617 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1234 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1233 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_155 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_620 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_619 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_618 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_617 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1232 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1231 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_616 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1232 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1231 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1230 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1229 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_615 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1230 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1229 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1228 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1227 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_614 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1228 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1227 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1226 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1225 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_613 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1226 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1225 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_154 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_616 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_615 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_614 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_613 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1224 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1223 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_612 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1224 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1223 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1222 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1221 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_611 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1222 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1221 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1220 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1219 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_610 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1220 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1219 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1218 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1217 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_609 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1218 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1217 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_153 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_612 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_611 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_610 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_609 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_39 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_156 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_155 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_154 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_153 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1216 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1215 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_608 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1216 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1215 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1214 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1213 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_607 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1214 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1213 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1212 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1211 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_606 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1212 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1211 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1210 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1209 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_605 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1210 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1209 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_152 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_608 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_607 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_606 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_605 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1208 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1207 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_604 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1208 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1207 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1206 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1205 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_603 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1206 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1205 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1204 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1203 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_602 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1204 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1203 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1202 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1201 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_601 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1202 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1201 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_151 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_604 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_603 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_602 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_601 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1200 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1199 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_600 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1200 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1199 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1198 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1197 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_599 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1198 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1197 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1196 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1195 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_598 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1196 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1195 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1194 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1193 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_597 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1194 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1193 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_150 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_600 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_599 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_598 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_597 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1192 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1191 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_596 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1192 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1191 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1190 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1189 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_595 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1190 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1189 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1188 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1187 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_594 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1188 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1187 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1186 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1185 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_593 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1186 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1185 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_149 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_596 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_595 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_594 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_593 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_38 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_152 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_151 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_150 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_149 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1184 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1183 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_592 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1184 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1183 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1182 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1181 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_591 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1182 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1181 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1180 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1179 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_590 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1180 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1179 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1178 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1177 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_589 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1178 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1177 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_148 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_592 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_591 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_590 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_589 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1176 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1175 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_588 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1176 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1175 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1174 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1173 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_587 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1174 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1173 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1172 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1171 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_586 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1172 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1171 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1170 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1169 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_585 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1170 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1169 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_147 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_588 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_587 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_586 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_585 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1168 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1167 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_584 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1168 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1167 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1166 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1165 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_583 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1166 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1165 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1164 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1163 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_582 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1164 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1163 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1162 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1161 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_581 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1162 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1161 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_146 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_584 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_583 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_582 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_581 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1160 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1159 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_580 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1160 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1159 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1158 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1157 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_579 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1158 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1157 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1156 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1155 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_578 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1156 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1155 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1154 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1153 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_577 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1154 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1153 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_145 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_580 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_579 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_578 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_577 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_37 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_148 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_147 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_146 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_145 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_10 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U6 ( .A(s84[3]), .B(n2), .C(s83[3]), .D(n1), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n2), .C(s83[2]), .D(n1), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n2), .C(s83[1]), .D(n1), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n2), .C(s83[0]), .D(n1), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n3), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n3), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n3), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n3), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n2), .C(c_out810), .D(n1), .Z(c_out8) );
  bit4_40 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_39 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_38 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_37 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVDX1 U3 ( .A(n5), .Z0(n2), .Z1(n1) );
  CANR2X1 U4 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n3), .Z(n5) );
  CIVX2 U5 ( .A(c_in8), .Z(n3) );
endmodule


module Add_half_1152 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1151 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_576 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1152 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1151 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1150 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1149 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_575 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1150 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1149 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1148 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1147 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_574 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1148 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1147 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1146 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1145 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_573 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1146 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1145 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_144 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n2), .Z(c_out2) );
  Add_full_576 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_575 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_574 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_573 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n3), .Z(n1) );
  CANR2XL U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n3), .Z(n2) );
  CAOR2XL U5 ( .A(s4), .B(n1), .C(s3), .D(n2), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_1144 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1143 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_572 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1144 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1143 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1142 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1141 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_571 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1142 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1141 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1140 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1139 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_570 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1140 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1139 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1138 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1137 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_569 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1138 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1137 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_143 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_572 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_571 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_570 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_569 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1136 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1135 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_568 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1136 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1135 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1134 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1133 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_567 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1134 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1133 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1132 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1131 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_566 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1132 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1131 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1130 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1129 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_565 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1130 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1129 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_142 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_568 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_567 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_566 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_565 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1128 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1127 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_564 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1128 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1127 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1126 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1125 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_563 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1126 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1125 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1124 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1123 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_562 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1124 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1123 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1122 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1121 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_561 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1122 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1121 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_141 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_564 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_563 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_562 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_561 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U5 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_36 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_144 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_143 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_142 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_141 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(n2), .D(c_out400), .Z(n3) );
  CAOR2XL U4 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1120 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1119 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_560 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1120 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1119 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1118 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1117 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_559 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1118 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1117 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1116 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1115 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_558 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1116 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1115 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1114 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1113 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_557 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1114 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1113 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_140 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_560 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_559 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_558 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_557 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1112 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1111 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_556 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1112 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1111 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1110 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1109 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_555 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1110 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1109 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1108 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1107 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_554 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1108 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1107 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1106 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1105 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_553 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1106 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1105 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_139 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_556 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_555 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_554 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_553 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1104 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1103 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_552 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1104 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1103 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1102 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1101 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_551 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1102 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1101 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1100 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1099 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_550 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1100 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1099 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1098 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1097 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_549 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1098 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1097 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_138 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  Add_full_552 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_551 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_550 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_549 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U8 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1096 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1095 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_548 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1096 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1095 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1094 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1093 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_547 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1094 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1093 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1092 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1091 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_546 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1092 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1091 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1090 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1089 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_545 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1090 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1089 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_137 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_548 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_547 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_546 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_545 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_35 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_140 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_139 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_138 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_137 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1088 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1087 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_544 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1088 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1087 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1086 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1085 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_543 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1086 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1085 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1084 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1083 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_542 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1084 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1083 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1082 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1081 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_541 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1082 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1081 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_136 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_544 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_543 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_542 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_541 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1080 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1079 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_540 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1080 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1079 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1078 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1077 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_539 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1078 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1077 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1076 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1075 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_538 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1076 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1075 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1074 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1073 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_537 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1074 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1073 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_135 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_540 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_539 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_538 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_537 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1072 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1071 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_536 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1072 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1071 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1070 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1069 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_535 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1070 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1069 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1068 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1067 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_534 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1068 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1067 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1066 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1065 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_533 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1066 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1065 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_134 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_536 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_535 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_534 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_533 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1064 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1063 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_532 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1064 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1063 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1062 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1061 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_531 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1062 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1061 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1060 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1059 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_530 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1060 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1059 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1058 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1057 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_529 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1058 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1057 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_133 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_532 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_531 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_530 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_529 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_34 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_136 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_135 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_134 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_133 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_1056 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1055 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_528 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1056 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1055 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1054 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1053 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_527 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1054 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1053 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1052 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1051 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_526 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1052 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1051 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1050 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1049 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_525 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1050 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1049 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_132 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_528 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_527 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_526 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_525 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1048 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1047 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_524 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1048 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1047 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1046 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1045 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_523 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1046 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1045 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1044 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1043 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_522 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1044 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1043 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1042 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1041 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_521 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1042 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1041 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_131 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_524 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_523 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_522 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_521 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1040 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1039 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_520 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1040 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1039 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1038 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1037 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_519 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1038 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1037 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1036 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1035 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_518 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1036 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1035 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1034 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1033 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_517 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1034 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1033 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_130 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_520 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_519 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_518 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_517 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1032 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1031 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_516 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1032 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1031 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1030 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1029 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_515 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1030 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1029 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1028 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1027 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_514 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1028 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1027 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1026 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1025 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_513 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1026 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1025 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_129 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_516 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_515 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_514 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_513 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_33 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_132 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_131 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_130 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_129 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_9 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U6 ( .A(s84[3]), .B(n1), .C(s83[3]), .D(n3), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n1), .C(s83[2]), .D(n3), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n1), .C(s83[1]), .D(n3), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n1), .C(s83[0]), .D(n3), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n2), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n2), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n2), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n2), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n1), .C(c_out810), .D(n3), .Z(c_out8) );
  bit4_36 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_35 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_34 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_33 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CANR2X2 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in8), .Z(n2) );
endmodule


module bit16_3 ( sum16, c_out16, a16, b16, c_in16 );
  output [15:0] sum16;
  input [15:0] a16;
  input [15:0] b16;
  input c_in16;
  output c_out16;
  wire   c_out1600, c_out1601, c_out1610, c_out1611, n1, n2, n3, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36;
  wire   [7:0] s161;
  wire   [7:0] s162;
  wire   [7:0] s163;
  wire   [7:0] s164;

  CAOR2X1 U8 ( .A(s162[7]), .B(c_in16), .C(s161[7]), .D(n35), .Z(sum16[7]) );
  CAOR2X1 U9 ( .A(s162[6]), .B(c_in16), .C(s161[6]), .D(n35), .Z(sum16[6]) );
  CAOR2X1 U10 ( .A(s162[5]), .B(c_in16), .C(s161[5]), .D(n35), .Z(sum16[5]) );
  CAOR2X1 U11 ( .A(s162[4]), .B(c_in16), .C(s161[4]), .D(n35), .Z(sum16[4]) );
  CAOR2X1 U12 ( .A(s162[3]), .B(c_in16), .C(s161[3]), .D(n35), .Z(sum16[3]) );
  CAOR2X1 U13 ( .A(s162[2]), .B(c_in16), .C(s161[2]), .D(n35), .Z(sum16[2]) );
  CAOR2X1 U14 ( .A(s162[1]), .B(c_in16), .C(s161[1]), .D(n35), .Z(sum16[1]) );
  CAOR2X1 U21 ( .A(s162[0]), .B(c_in16), .C(s161[0]), .D(n35), .Z(sum16[0]) );
  bit8_12 A161 ( .sum8(s161), .c_out8(c_out1600), .a8({n26, n25, n24, n6, n23, 
        n22, n5, n21}), .b8({n13, n1, n12, n11, n2, n10, n9, n8}), .c_in8(1'b0) );
  bit8_11 A162 ( .sum8(s162), .c_out8(c_out1601), .a8({n26, n25, n24, n6, n23, 
        n22, n5, n21}), .b8({n13, n1, n12, n11, n2, n10, n9, n8}), .c_in8(1'b1) );
  bit8_10 A163 ( .sum8(s163), .c_out8(c_out1610), .a8({n33, n32, n31, n30, n29, 
        n28, n27, n7}), .b8({n20, n19, b16[13], n18, n17, n16, n15, n14}), 
        .c_in8(1'b0) );
  bit8_9 A164 ( .sum8(s164), .c_out8(c_out1611), .a8({n33, n32, n31, n30, n29, 
        n28, n27, n7}), .b8({n20, n19, b16[13], n18, n17, n16, n15, n14}), 
        .c_in8(1'b1) );
  CNIVX3 U3 ( .A(a16[8]), .Z(n7) );
  CNIVX2 U4 ( .A(b16[3]), .Z(n2) );
  CNIVX2 U5 ( .A(b16[6]), .Z(n1) );
  CNIVX1 U6 ( .A(b16[5]), .Z(n12) );
  CNIVX2 U7 ( .A(a16[1]), .Z(n5) );
  CNIVX16 U15 ( .A(a16[0]), .Z(n21) );
  CNIVX2 U16 ( .A(a16[2]), .Z(n22) );
  CNIVX2 U17 ( .A(a16[4]), .Z(n6) );
  CIVX2 U18 ( .A(n36), .Z(n34) );
  CIVXL U19 ( .A(n34), .Z(n3) );
  CANR2X2 U20 ( .A(c_out1601), .B(c_in16), .C(c_out1600), .D(n35), .Z(n36) );
  CNIVX2 U22 ( .A(a16[12]), .Z(n30) );
  CNIVX16 U23 ( .A(b16[0]), .Z(n8) );
  CNIVX2 U24 ( .A(a16[9]), .Z(n27) );
  CNIVX2 U25 ( .A(a16[6]), .Z(n25) );
  CNIVX2 U26 ( .A(a16[10]), .Z(n28) );
  CNIVX2 U27 ( .A(a16[3]), .Z(n23) );
  CNIVX2 U28 ( .A(a16[5]), .Z(n24) );
  CNIVX2 U29 ( .A(b16[2]), .Z(n10) );
  CNIVX2 U30 ( .A(b16[4]), .Z(n11) );
  CAOR2X1 U31 ( .A(c_out1611), .B(n34), .C(c_out1610), .D(n36), .Z(c_out16) );
  CNIVX1 U32 ( .A(a16[13]), .Z(n31) );
  CNIVX1 U33 ( .A(b16[15]), .Z(n20) );
  CNIVX1 U34 ( .A(b16[14]), .Z(n19) );
  CNIVX1 U35 ( .A(b16[11]), .Z(n17) );
  CNIVX1 U36 ( .A(b16[7]), .Z(n13) );
  CNIVX1 U37 ( .A(a16[15]), .Z(n33) );
  CNIVX1 U38 ( .A(a16[11]), .Z(n29) );
  CNIVX1 U39 ( .A(a16[7]), .Z(n26) );
  CNIVX1 U40 ( .A(a16[14]), .Z(n32) );
  CNIVX2 U41 ( .A(b16[9]), .Z(n15) );
  CNIVX2 U42 ( .A(b16[10]), .Z(n16) );
  CNIVX2 U43 ( .A(b16[8]), .Z(n14) );
  CNIVX2 U44 ( .A(b16[1]), .Z(n9) );
  CAOR2XL U45 ( .A(s164[6]), .B(n34), .C(s163[6]), .D(n3), .Z(sum16[14]) );
  CAOR2XL U46 ( .A(s164[5]), .B(n34), .C(s163[5]), .D(n3), .Z(sum16[13]) );
  CAOR2XL U47 ( .A(s164[4]), .B(n34), .C(s163[4]), .D(n3), .Z(sum16[12]) );
  CAOR2XL U48 ( .A(s164[3]), .B(n34), .C(s163[3]), .D(n3), .Z(sum16[11]) );
  CAOR2XL U49 ( .A(s164[2]), .B(n34), .C(s163[2]), .D(n36), .Z(sum16[10]) );
  CNIVX2 U50 ( .A(b16[12]), .Z(n18) );
  CAOR2XL U51 ( .A(s164[1]), .B(n34), .C(s163[1]), .D(n3), .Z(sum16[9]) );
  CAOR2XL U52 ( .A(s164[0]), .B(n34), .C(s163[0]), .D(n3), .Z(sum16[8]) );
  CAOR2XL U53 ( .A(s164[7]), .B(n34), .C(s163[7]), .D(n3), .Z(sum16[15]) );
  CIVX2 U54 ( .A(c_in16), .Z(n35) );
endmodule


module Add_half_1024 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1023 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_512 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1024 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1023 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1022 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1021 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_511 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1022 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1021 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1020 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1019 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_510 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1020 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1019 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1018 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1017 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_509 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1018 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1017 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_128 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_512 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_511 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_510 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_509 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1016 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1015 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_508 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1016 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1015 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1014 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1013 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_507 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1014 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1013 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1012 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1011 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_506 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1012 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1011 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1010 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1009 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_505 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1010 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1009 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_127 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_508 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_507 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_506 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_505 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1008 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1007 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_504 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1008 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1007 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1006 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1005 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_503 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1006 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1005 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1004 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1003 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_502 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1004 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1003 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_1002 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1001 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_501 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1002 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1001 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_126 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_504 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_503 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_502 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_501 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_1000 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_999 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_500 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_1000 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_999 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_998 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_997 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_499 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_998 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_997 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_996 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_995 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_498 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_996 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_995 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_994 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_993 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_497 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_994 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_993 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_125 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_500 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_499 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_498 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_497 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_32 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_128 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_127 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_126 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_125 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2XL U5 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CIVX2 U6 ( .A(n3), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_992 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_991 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_496 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_992 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_991 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_990 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_989 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_495 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_990 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_989 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_988 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_987 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_494 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_988 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_987 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_986 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_985 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_493 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_986 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_985 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_124 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_496 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_495 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_494 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_493 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_984 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_983 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_492 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_984 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_983 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_982 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_981 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_491 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_982 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_981 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_980 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_979 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_490 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_980 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_979 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_978 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_977 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_489 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_978 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_977 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_123 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_492 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_491 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_490 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_489 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_976 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_975 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_488 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_976 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_975 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_974 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_973 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_487 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_974 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_973 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_972 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_971 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_486 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_972 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_971 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_970 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_969 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_485 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_970 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_969 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_122 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  Add_full_488 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_487 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_486 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_485 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U8 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_968 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_967 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_484 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_968 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_967 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_966 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_965 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_483 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_966 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_965 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_964 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_963 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_482 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_964 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_963 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_962 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_961 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_481 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_962 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_961 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_121 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_484 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_483 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_482 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_481 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_31 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_124 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_123 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_122 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_121 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_960 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_959 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_480 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_960 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_959 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_958 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_957 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_479 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_958 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_957 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_956 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_955 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_478 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_956 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_955 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_954 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_953 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_477 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_954 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_953 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_120 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_480 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_479 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_478 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_477 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_952 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_951 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_476 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_952 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_951 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_950 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_949 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_475 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_950 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_949 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_948 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_947 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_474 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_948 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_947 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_946 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_945 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_473 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_946 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_945 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_119 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_476 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_475 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_474 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_473 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_944 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_943 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_472 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_944 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_943 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_942 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_941 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_471 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_942 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_941 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_940 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_939 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_470 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_940 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_939 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_938 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_937 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_469 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_938 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_937 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_118 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_472 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_471 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_470 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_469 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_936 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_935 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_468 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_936 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_935 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_934 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_933 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_467 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_934 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_933 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_932 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_931 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_466 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_932 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_931 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_930 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_929 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_465 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_930 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_929 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_117 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_468 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_467 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_466 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_465 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_30 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_120 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_119 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_118 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_117 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_928 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_927 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_464 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_928 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_927 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_926 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_925 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_463 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_926 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_925 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_924 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_923 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_462 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_924 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_923 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_922 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_921 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_461 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_922 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_921 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_116 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_464 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_463 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_462 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_461 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_920 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_919 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_460 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_920 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_919 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_918 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_917 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_459 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_918 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_917 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_916 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_915 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_458 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_916 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_915 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_914 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_913 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_457 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_914 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_913 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_115 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_460 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_459 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_458 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_457 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_912 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_911 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_456 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_912 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_911 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_910 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_909 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_455 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_910 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_909 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_908 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_907 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_454 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_908 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_907 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_906 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_905 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_453 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_906 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_905 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_114 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_456 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_455 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_454 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_453 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_904 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_903 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_452 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_904 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_903 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_902 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_901 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_451 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_902 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_901 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_900 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_899 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_450 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_900 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_899 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_898 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_897 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_449 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_898 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_897 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_113 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_452 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_451 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_450 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_449 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_29 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_116 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_115 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_114 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_113 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2XL U5 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CIVX2 U6 ( .A(n3), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_8 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n2), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n2), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n2), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n2), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n1), .C(c_out810), .D(n3), .Z(c_out8) );
  bit4_32 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_31 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_30 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_29 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CANR2X2 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s84[0]), .B(n1), .C(s83[0]), .D(n3), .Z(sum8[4]) );
  CAOR2XL U5 ( .A(s84[1]), .B(n1), .C(s83[1]), .D(n3), .Z(sum8[5]) );
  CAOR2XL U6 ( .A(s84[2]), .B(n1), .C(s83[2]), .D(n3), .Z(sum8[6]) );
  CAOR2XL U7 ( .A(s84[3]), .B(n1), .C(s83[3]), .D(n3), .Z(sum8[7]) );
  CIVX2 U8 ( .A(n3), .Z(n1) );
  CIVX2 U9 ( .A(c_in8), .Z(n2) );
endmodule


module Add_half_896 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_895 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_448 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_896 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_895 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_894 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_893 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_447 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_894 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_893 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_892 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_891 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_446 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_892 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_891 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_890 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_889 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_445 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_890 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_889 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_112 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_448 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_447 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_446 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_445 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_888 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_887 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_444 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_888 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_887 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_886 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_885 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_443 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_886 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_885 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_884 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_883 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_442 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_884 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_883 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_882 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_881 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_441 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_882 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_881 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_111 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_444 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_443 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_442 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_441 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_880 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_879 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_440 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_880 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_879 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_878 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_877 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_439 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_878 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_877 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_876 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_875 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_438 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_876 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_875 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_874 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_873 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_437 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_874 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_873 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_110 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_440 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_439 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_438 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_437 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_872 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_871 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_436 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_872 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_871 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_870 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_869 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_435 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_870 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_869 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_868 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_867 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_434 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_868 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_867 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_866 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_865 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_433 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_866 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_865 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_109 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_436 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_435 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_434 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_433 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_28 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_112 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_111 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_110 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_109 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_864 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_863 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_432 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_864 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_863 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_862 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_861 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_431 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_862 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_861 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_860 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_859 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_430 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_860 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_859 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_858 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_857 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_429 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_858 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_857 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_108 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_432 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_431 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_430 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_429 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_856 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_855 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_428 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_856 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_855 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_854 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_853 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_427 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_854 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_853 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_852 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_851 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_426 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_852 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_851 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_850 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_849 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_425 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_850 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_849 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_107 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_428 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_427 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_426 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_425 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_848 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_847 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_424 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_848 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_847 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_846 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_845 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_423 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_846 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_845 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_844 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_843 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_422 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_844 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_843 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_842 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_841 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_421 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_842 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_841 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_106 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_424 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_423 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_422 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_421 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_840 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_839 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_420 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_840 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_839 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_838 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_837 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_419 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_838 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_837 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_836 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_835 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_418 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_836 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_835 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_834 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_833 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_417 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_834 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_833 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_105 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_420 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_419 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_418 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_417 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_27 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_108 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_107 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_106 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_105 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_832 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_831 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_416 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_832 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_831 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_830 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_829 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_415 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_830 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_829 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_828 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_827 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_414 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_828 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_827 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_826 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_825 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_413 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_826 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_825 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_104 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_416 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_415 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_414 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_413 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_824 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_823 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_412 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_824 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_823 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_822 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_821 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_411 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_822 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_821 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_820 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_819 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_410 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_820 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_819 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_818 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_817 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_409 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_818 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_817 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_103 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_412 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_411 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_410 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_409 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_816 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_815 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_408 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_816 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_815 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_814 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_813 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_407 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_814 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_813 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_812 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_811 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_406 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_812 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_811 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_810 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_809 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_405 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_810 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_809 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_102 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_408 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_407 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_406 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_405 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_808 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_807 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_404 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_808 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_807 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_806 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_805 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_403 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_806 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_805 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_804 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_803 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_402 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_804 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_803 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_802 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_801 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_401 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_802 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_801 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_101 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_404 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_403 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_402 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_401 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_26 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_104 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_103 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_102 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_101 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_800 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_799 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_400 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_800 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_799 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_798 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_797 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_399 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_798 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_797 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_796 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_795 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_398 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_796 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_795 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_794 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_793 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_397 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_794 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_793 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_100 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_400 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_399 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_398 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_397 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_792 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_791 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_396 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_792 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_791 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_790 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_789 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_395 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_790 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_789 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_788 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_787 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_394 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_788 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_787 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_786 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_785 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_393 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_786 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_785 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_99 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_396 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_395 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_394 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_393 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_784 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_783 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_392 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_784 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_783 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_782 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_781 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_391 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_782 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_781 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_780 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_779 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_390 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_780 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_779 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_778 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_777 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_389 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_778 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_777 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_98 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_392 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_391 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_390 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_389 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_776 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_775 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_388 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_776 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_775 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_774 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_773 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_387 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_774 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_773 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_772 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_771 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_386 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_772 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_771 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_770 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_769 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_385 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_770 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_769 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_97 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_388 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_387 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_386 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_385 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_25 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_100 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_99 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_98 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_97 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_7 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CANR2X2 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n2), .Z(n3) );
  CAOR2X1 U6 ( .A(s84[3]), .B(n1), .C(s83[3]), .D(n3), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n1), .C(s83[2]), .D(n3), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n1), .C(s83[1]), .D(n3), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n1), .C(s83[0]), .D(n3), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n2), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n2), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n2), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n2), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n1), .C(c_out810), .D(n3), .Z(c_out8) );
  bit4_28 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_27 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_26 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_25 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in8), .Z(n2) );
endmodule


module Add_half_768 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_767 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_384 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_768 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_767 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_766 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_765 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_383 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_766 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_765 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_764 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_763 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_382 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_764 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_763 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_762 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_761 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_381 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_762 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_761 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_96 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_384 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_383 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_382 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_381 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_760 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_759 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_380 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_760 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_759 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_758 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_757 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_379 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_758 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_757 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_756 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_755 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_378 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_756 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_755 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_754 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_753 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_377 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_754 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_753 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_95 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_380 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_379 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_378 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_377 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_752 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_751 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_376 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_752 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_751 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_750 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_749 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_375 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_750 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_749 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_748 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_747 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_374 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_748 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_747 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_746 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_745 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_373 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_746 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_745 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_94 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_376 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_375 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_374 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_373 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_744 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_743 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_372 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_744 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_743 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_742 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_741 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_371 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_742 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_741 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_740 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_739 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_370 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_740 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_739 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_738 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_737 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_369 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_738 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_737 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_93 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_372 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_371 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_370 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_369 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_24 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_96 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_95 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_94 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_93 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_736 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_735 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_368 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_736 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_735 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_734 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_733 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_367 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_734 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_733 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_732 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_731 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_366 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_732 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_731 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_730 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_729 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_365 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_730 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_729 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_92 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_368 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_367 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_366 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_365 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_728 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_727 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_364 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_728 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_727 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_726 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_725 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_363 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_726 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_725 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_724 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_723 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_362 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_724 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_723 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_722 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_721 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_361 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_722 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_721 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_91 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_364 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_363 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_362 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_361 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_720 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_719 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_360 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_720 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_719 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_718 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_717 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_359 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_718 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_717 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_716 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_715 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_358 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_716 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_715 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_714 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_713 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_357 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_714 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_713 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_90 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_360 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_359 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_358 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_357 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_712 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_711 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_356 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_712 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_711 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_710 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_709 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_355 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_710 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_709 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_708 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_707 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_354 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_708 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_707 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_706 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_705 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_353 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_706 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_705 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_89 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_356 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_355 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_354 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_353 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_23 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_92 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_91 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_90 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_89 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_704 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_703 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_352 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_704 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_703 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_702 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_701 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_351 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_702 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_701 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_700 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_699 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_350 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_700 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_699 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_698 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_697 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_349 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_698 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_697 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_88 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_352 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_351 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_350 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_349 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_696 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_695 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_348 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_696 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_695 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_694 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_693 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_347 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_694 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_693 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_692 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_691 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_346 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_692 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_691 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_690 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_689 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_345 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_690 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_689 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_87 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_348 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_347 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_346 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_345 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_688 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_687 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_344 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_688 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_687 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_686 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_685 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_343 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_686 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_685 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_684 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_683 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_342 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_684 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_683 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_682 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_681 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_341 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_682 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_681 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_86 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_344 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_343 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_342 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_341 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_680 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_679 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_340 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_680 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_679 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_678 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_677 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_339 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_678 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_677 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_676 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_675 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_338 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_676 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_675 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_674 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_673 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_337 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_674 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_673 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_85 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_340 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_339 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_338 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_337 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_22 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_88 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_87 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_86 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_85 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_672 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_671 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_336 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_672 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_671 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_670 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_669 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_335 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_670 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_669 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_668 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_667 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_334 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_668 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_667 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_666 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_665 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_333 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_666 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_665 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_84 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_336 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_335 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_334 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_333 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_664 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_663 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_332 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_664 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_663 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_662 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_661 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_331 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_662 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_661 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_660 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_659 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_330 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_660 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_659 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_658 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_657 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_329 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_658 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_657 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_83 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_332 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_331 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_330 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_329 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_656 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_655 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_328 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_656 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_655 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_654 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_653 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_327 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_654 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_653 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_652 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_651 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_326 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_652 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_651 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_650 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_649 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_325 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_650 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_649 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_82 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_328 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_327 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_326 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_325 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_648 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_647 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_324 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_648 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_647 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_646 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_645 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_323 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_646 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_645 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_644 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_643 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_322 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_644 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_643 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_642 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_641 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_321 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_642 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_641 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_81 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_324 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_323 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_322 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_321 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_21 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_84 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_83 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_82 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_81 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_6 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U6 ( .A(s84[3]), .B(n1), .C(s83[3]), .D(n3), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n1), .C(s83[2]), .D(n3), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n1), .C(s83[1]), .D(n3), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n1), .C(s83[0]), .D(n3), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n2), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n2), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n2), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n2), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n1), .C(c_out810), .D(n3), .Z(c_out8) );
  bit4_24 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_23 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_22 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_21 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CANR2X1 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in8), .Z(n2) );
endmodule


module Add_half_640 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_639 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_320 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_640 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_639 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_638 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_637 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_319 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_638 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_637 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_636 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_635 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_318 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_636 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_635 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_634 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_633 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_317 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_634 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_633 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_80 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_320 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_319 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_318 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_317 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_632 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_631 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_316 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_632 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_631 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_630 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_629 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_315 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_630 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_629 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_628 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_627 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_314 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_628 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_627 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_626 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_625 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_313 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_626 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_625 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_79 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_316 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_315 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_314 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_313 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_624 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_623 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_312 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_624 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_623 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_622 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_621 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_311 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_622 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_621 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_620 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_619 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_310 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_620 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_619 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_618 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_617 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_309 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_618 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_617 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_78 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_312 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_311 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_310 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_309 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_616 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_615 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_308 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_616 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_615 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_614 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_613 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_307 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_614 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_613 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_612 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_611 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_306 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_612 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_611 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_610 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_609 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_305 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_610 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_609 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_77 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_308 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_307 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_306 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_305 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_20 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_80 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_79 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_78 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_77 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_608 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_607 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_304 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_608 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_607 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_606 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_605 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_303 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_606 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_605 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_604 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_603 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_302 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_604 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_603 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_602 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_601 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_301 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_602 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_601 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_76 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_304 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_303 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_302 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_301 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_600 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_599 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_300 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_600 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_599 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_598 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_597 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_299 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_598 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_597 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_596 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_595 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_298 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_596 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_595 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_594 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_593 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_297 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_594 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_593 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_75 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_300 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_299 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_298 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_297 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_592 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_591 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_296 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_592 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_591 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_590 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_589 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_295 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_590 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_589 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_588 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_587 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_294 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_588 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_587 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_586 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_585 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_293 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_586 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_585 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_74 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_296 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_295 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_294 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_293 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_584 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_583 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_292 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_584 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_583 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_582 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_581 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_291 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_582 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_581 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_580 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_579 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_290 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_580 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_579 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_578 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_577 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_289 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_578 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_577 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_73 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_292 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_291 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_290 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_289 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_19 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_76 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_75 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_74 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_73 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_576 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_575 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_288 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_576 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_575 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_574 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_573 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_287 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_574 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_573 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_572 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_571 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_286 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_572 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_571 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_570 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_569 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_285 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_570 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_569 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_72 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_288 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_287 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_286 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_285 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_568 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_567 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_284 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_568 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_567 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_566 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_565 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_283 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_566 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_565 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_564 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_563 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_282 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_564 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_563 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_562 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_561 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_281 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_562 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_561 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_71 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_284 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_283 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_282 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_281 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_560 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_559 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_280 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_560 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_559 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_558 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_557 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_279 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_558 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_557 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_556 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_555 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_278 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_556 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_555 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_554 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_553 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_277 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_554 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_553 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_70 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_280 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_279 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_278 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_277 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_552 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_551 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_276 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_552 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_551 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_550 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_549 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_275 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_550 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_549 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_548 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_547 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_274 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_548 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_547 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_546 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_545 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_273 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_546 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_545 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_69 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_276 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_275 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_274 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_273 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_18 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_72 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_71 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_70 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_69 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_544 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_543 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_272 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_544 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_543 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_542 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_541 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_271 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_542 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_541 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_540 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_539 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_270 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_540 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_539 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_538 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_537 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_269 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_538 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_537 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_68 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_272 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_271 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_270 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_269 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_536 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_535 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_268 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_536 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_535 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_534 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_533 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_267 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_534 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_533 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_532 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_531 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_266 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_532 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_531 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_530 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_529 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_265 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_530 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_529 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_67 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_268 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_267 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_266 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_265 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_528 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_527 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_264 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_528 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_527 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_526 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_525 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_263 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_526 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_525 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_524 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_523 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_262 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_524 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_523 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_522 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_521 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_261 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_522 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_521 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_66 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_264 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_263 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_262 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_261 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_520 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_519 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_260 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_520 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_519 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_518 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_517 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_259 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_518 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_517 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_516 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_515 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_258 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_516 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_515 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_514 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_513 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_257 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_514 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_513 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_65 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_260 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_259 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_258 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_257 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_17 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_68 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_67 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_66 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_65 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_5 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U6 ( .A(s84[3]), .B(n1), .C(s83[3]), .D(n3), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n1), .C(s83[2]), .D(n3), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n1), .C(s83[1]), .D(n3), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n1), .C(s83[0]), .D(n3), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n2), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n2), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n2), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n2), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n1), .C(c_out810), .D(n3), .Z(c_out8) );
  bit4_20 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_19 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_18 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_17 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CANR2X1 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in8), .Z(n2) );
endmodule


module bit16_2 ( sum16, c_out16, a16, b16, c_in16 );
  output [15:0] sum16;
  input [15:0] a16;
  input [15:0] b16;
  input c_in16;
  output c_out16;
  wire   c_out1600, c_out1601, c_out1610, c_out1611, n1, n2, n3, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37;
  wire   [7:0] s161;
  wire   [7:0] s162;
  wire   [7:0] s163;
  wire   [7:0] s164;

  CAOR2X1 U6 ( .A(s164[1]), .B(n3), .C(s163[1]), .D(n2), .Z(sum16[9]) );
  CAOR2X1 U7 ( .A(s164[0]), .B(n3), .C(s163[0]), .D(n2), .Z(sum16[8]) );
  CAOR2X1 U8 ( .A(s162[7]), .B(c_in16), .C(s161[7]), .D(n36), .Z(sum16[7]) );
  CAOR2X1 U9 ( .A(s162[6]), .B(c_in16), .C(s161[6]), .D(n36), .Z(sum16[6]) );
  CAOR2X1 U10 ( .A(s162[5]), .B(c_in16), .C(s161[5]), .D(n36), .Z(sum16[5]) );
  CAOR2X1 U11 ( .A(s162[4]), .B(c_in16), .C(s161[4]), .D(n36), .Z(sum16[4]) );
  CAOR2X1 U12 ( .A(s162[3]), .B(c_in16), .C(s161[3]), .D(n36), .Z(sum16[3]) );
  CAOR2X1 U13 ( .A(s162[2]), .B(c_in16), .C(s161[2]), .D(n36), .Z(sum16[2]) );
  CAOR2X1 U14 ( .A(s162[1]), .B(c_in16), .C(s161[1]), .D(n36), .Z(sum16[1]) );
  CAOR2X1 U15 ( .A(s164[7]), .B(n3), .C(s163[7]), .D(n2), .Z(sum16[15]) );
  CAOR2X1 U16 ( .A(s164[6]), .B(n3), .C(s163[6]), .D(n2), .Z(sum16[14]) );
  CAOR2X1 U17 ( .A(s164[5]), .B(n3), .C(s163[5]), .D(n2), .Z(sum16[13]) );
  CAOR2X1 U18 ( .A(s164[4]), .B(n3), .C(s163[4]), .D(n2), .Z(sum16[12]) );
  CAOR2X1 U19 ( .A(s164[3]), .B(n3), .C(s163[3]), .D(n2), .Z(sum16[11]) );
  CAOR2X1 U20 ( .A(s164[2]), .B(n3), .C(s163[2]), .D(n2), .Z(sum16[10]) );
  CAOR2X1 U21 ( .A(s162[0]), .B(c_in16), .C(s161[0]), .D(n36), .Z(sum16[0]) );
  CAOR2X1 U22 ( .A(c_out1611), .B(n3), .C(c_out1610), .D(n2), .Z(c_out16) );
  bit8_8 A161 ( .sum8(s161), .c_out8(c_out1600), .a8({n27, n26, n25, n1, n24, 
        n23, n22, n5}), .b8({n13, n12, n11, n10, n9, n8, n7, n6}), .c_in8(1'b0) );
  bit8_7 A162 ( .sum8(s162), .c_out8(c_out1601), .a8({n27, n26, n25, n1, n24, 
        n23, n22, n5}), .b8({n13, n12, n11, n10, n9, n8, n7, n6}), .c_in8(1'b1) );
  bit8_6 A163 ( .sum8(s163), .c_out8(c_out1610), .a8({n35, n34, n33, n32, n31, 
        n30, n29, n28}), .b8({n21, n20, n19, n18, n17, n16, n15, n14}), 
        .c_in8(1'b0) );
  bit8_5 A164 ( .sum8(s164), .c_out8(c_out1611), .a8({n35, n34, n33, n32, n31, 
        n30, n29, n28}), .b8({n21, n20, n19, n18, n17, n16, n15, n14}), 
        .c_in8(1'b1) );
  CNIVX2 U3 ( .A(a16[4]), .Z(n1) );
  CNIVX2 U4 ( .A(b16[2]), .Z(n8) );
  CNIVX2 U5 ( .A(b16[4]), .Z(n10) );
  CNIVX2 U23 ( .A(b16[1]), .Z(n7) );
  CNIVX2 U24 ( .A(a16[0]), .Z(n5) );
  CNIVX1 U25 ( .A(b16[8]), .Z(n14) );
  CIVDX1 U26 ( .A(n37), .Z0(n3), .Z1(n2) );
  CANR2X1 U27 ( .A(c_out1601), .B(c_in16), .C(c_out1600), .D(n36), .Z(n37) );
  CNIVX2 U28 ( .A(b16[0]), .Z(n6) );
  CNIVX1 U29 ( .A(a16[8]), .Z(n28) );
  CNIVX1 U30 ( .A(a16[2]), .Z(n23) );
  CNIVX1 U31 ( .A(a16[1]), .Z(n22) );
  CNIVX1 U32 ( .A(b16[6]), .Z(n12) );
  CNIVX1 U33 ( .A(b16[5]), .Z(n11) );
  CNIVX1 U34 ( .A(b16[10]), .Z(n16) );
  CNIVX1 U35 ( .A(b16[9]), .Z(n15) );
  CNIVX1 U36 ( .A(b16[11]), .Z(n17) );
  CNIVX1 U37 ( .A(b16[13]), .Z(n19) );
  CNIVX1 U38 ( .A(b16[14]), .Z(n20) );
  CNIVX1 U39 ( .A(b16[7]), .Z(n13) );
  CNIVX1 U40 ( .A(b16[3]), .Z(n9) );
  CNIVX1 U41 ( .A(b16[12]), .Z(n18) );
  CNIVX1 U42 ( .A(b16[15]), .Z(n21) );
  CNIVX1 U43 ( .A(a16[12]), .Z(n32) );
  CNIVX1 U44 ( .A(a16[11]), .Z(n31) );
  CNIVX1 U45 ( .A(a16[13]), .Z(n33) );
  CNIVX1 U46 ( .A(a16[14]), .Z(n34) );
  CNIVX1 U47 ( .A(a16[7]), .Z(n27) );
  CNIVX1 U48 ( .A(a16[15]), .Z(n35) );
  CNIVX1 U49 ( .A(a16[9]), .Z(n29) );
  CNIVX1 U50 ( .A(a16[3]), .Z(n24) );
  CNIVX1 U51 ( .A(a16[5]), .Z(n25) );
  CNIVX1 U52 ( .A(a16[6]), .Z(n26) );
  CNIVX1 U53 ( .A(a16[10]), .Z(n30) );
  CIVX2 U54 ( .A(c_in16), .Z(n36) );
endmodule


module Add_half_512 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_511 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_256 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_512 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_511 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_510 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_509 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_255 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_510 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_509 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_508 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_507 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_254 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_508 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_507 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_506 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_505 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_253 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_506 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_505 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_64 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_256 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_255 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_254 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_253 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_504 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(a), .Z(n1) );
  CENX1 U2 ( .A(b), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_503 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_252 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_504 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_503 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_502 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_501 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_251 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_502 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_501 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_500 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_499 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_250 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_500 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_499 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_498 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_497 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_249 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_498 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_497 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_63 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_252 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_251 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_250 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_249 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_496 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_495 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_248 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_496 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_495 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_494 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_493 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_247 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_494 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_493 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_492 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_491 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_246 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_492 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_491 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_490 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_489 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_245 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_490 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_489 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_62 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_248 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_247 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_246 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_245 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_488 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_487 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_244 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_488 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_487 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_486 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_485 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_243 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_486 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_485 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_484 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_483 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_242 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_484 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_483 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_482 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_481 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_241 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_482 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_481 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_61 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_244 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_243 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_242 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_241 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_16 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_64 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_63 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_62 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_61 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2XL U5 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CIVX2 U6 ( .A(n3), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_480 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_479 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_240 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_480 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_479 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_478 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_477 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_239 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_478 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_477 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_476 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_475 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_238 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_476 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_475 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_474 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_473 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_237 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_474 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_473 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_60 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_240 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_239 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_238 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_237 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_472 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_471 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_236 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_472 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_471 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_470 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_469 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_235 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_470 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_469 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_468 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_467 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_234 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_468 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_467 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_466 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_465 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_233 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_466 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_465 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_59 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_236 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_235 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_234 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_233 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_464 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_463 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_232 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_464 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_463 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_462 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_461 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_231 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_462 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_461 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_460 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_459 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_230 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_460 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_459 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_458 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_457 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_229 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_458 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_457 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_58 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_232 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_231 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_230 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_229 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_456 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_455 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_228 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_456 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_455 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_454 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_453 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_227 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_454 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_453 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_452 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_451 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_226 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_452 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_451 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_450 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_449 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_225 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_450 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_449 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_57 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_228 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_227 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_226 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_225 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_15 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_60 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_59 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_58 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_57 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_448 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_447 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_224 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_448 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_447 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_446 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_445 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_223 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_446 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_445 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_444 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_443 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_222 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_444 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_443 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_442 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_441 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_221 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_442 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_441 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_56 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_224 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_223 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_222 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_221 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_440 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_439 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_220 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_440 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_439 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_438 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_437 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_219 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_438 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_437 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_436 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_435 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_218 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_436 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_435 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_434 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_433 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_217 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_434 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_433 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_55 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_220 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_219 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_218 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_217 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_432 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_431 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_216 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_432 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_431 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_430 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_429 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_215 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_430 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_429 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_428 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_427 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_214 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_428 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_427 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_426 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_425 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_213 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_426 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_425 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_54 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_216 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_215 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_214 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_213 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_424 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_423 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_212 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_424 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_423 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_422 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_421 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_211 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_422 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_421 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_420 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_419 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_210 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_420 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_419 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_418 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_417 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_209 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_418 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_417 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_53 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_212 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_211 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_210 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_209 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_14 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_56 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_55 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_54 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_53 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2XL U3 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CIVX1 U4 ( .A(n3), .Z(n1) );
  CANR2X1 U5 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_416 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_415 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_208 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_416 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_415 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_414 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_413 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_207 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_414 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_413 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_412 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_411 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_206 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_412 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_411 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_410 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_409 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_205 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_410 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_409 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_52 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_208 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_207 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_206 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_205 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_408 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(a), .Z(n1) );
  CENX1 U2 ( .A(b), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_407 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_204 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_408 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_407 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_406 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_405 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_203 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_406 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_405 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_404 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_403 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_202 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_404 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_403 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_402 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_401 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_201 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_402 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_401 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_51 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_204 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_203 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_202 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_201 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_400 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_399 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_200 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_400 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_399 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_398 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_397 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_199 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_398 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_397 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_396 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_395 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_198 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_396 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_395 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_394 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_393 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_197 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_394 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_393 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_50 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_200 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_199 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_198 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_197 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_392 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_391 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_196 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_392 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_391 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_390 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_389 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_195 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_390 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_389 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_388 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_387 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_194 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_388 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_387 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_386 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_385 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_193 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_386 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_385 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_49 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_196 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_195 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_194 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_193 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_13 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n3), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n3), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n2), .Z(c_out4) );
  bit2_52 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_51 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_50 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_49 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n3), .Z(n1) );
  CIVXL U4 ( .A(n1), .Z(n2) );
  CAOR2XL U5 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n2), .Z(sum4[2]) );
  CAOR2XL U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n2), .Z(sum4[3]) );
  CIVX2 U7 ( .A(c_in4), .Z(n3) );
endmodule


module bit8_4 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n3), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n3), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n3), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n3), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n1), .C(c_out810), .D(n2), .Z(c_out8) );
  bit4_16 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_15 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_14 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_13 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVDX1 U3 ( .A(n5), .Z0(n1), .Z1(n2) );
  CANR2X1 U4 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n3), .Z(n5) );
  CAOR2XL U5 ( .A(s84[0]), .B(n1), .C(s83[0]), .D(n2), .Z(sum8[4]) );
  CAOR2XL U6 ( .A(s84[1]), .B(n1), .C(s83[1]), .D(n2), .Z(sum8[5]) );
  CAOR2XL U7 ( .A(s84[3]), .B(n1), .C(s83[3]), .D(n2), .Z(sum8[7]) );
  CAOR2XL U8 ( .A(s84[2]), .B(n1), .C(s83[2]), .D(n2), .Z(sum8[6]) );
  CIVX2 U9 ( .A(c_in8), .Z(n3) );
endmodule


module Add_half_384 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_383 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_192 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_384 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_383 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_382 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_381 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_191 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_382 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_381 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_380 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_379 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_190 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_380 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_379 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_378 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_377 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_189 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_378 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_377 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_48 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_192 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_191 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_190 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_189 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_376 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_375 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_188 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_376 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_375 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_374 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_373 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_187 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_374 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_373 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_372 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_371 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_186 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_372 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_371 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_370 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_369 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_185 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_370 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_369 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_47 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_188 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_187 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_186 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_185 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_368 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_367 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_184 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_368 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_367 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_366 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_365 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_183 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_366 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_365 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_364 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_363 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_182 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_364 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_363 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_362 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_361 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_181 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_362 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_361 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_46 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_184 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_183 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_182 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_181 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_360 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_359 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_180 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_360 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_359 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_358 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_357 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_179 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_358 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_357 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_356 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_355 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_178 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_356 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_355 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_354 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_353 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_177 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_354 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_353 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_45 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_180 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_179 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_178 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_177 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_12 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_48 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_47 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_46 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_45 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CAOR2XL U4 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2XL U5 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CIVX2 U6 ( .A(n3), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_352 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_351 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_176 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_352 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_351 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_350 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_349 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_175 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_350 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_349 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_348 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_347 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_174 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_348 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_347 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_346 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_345 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_173 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_346 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_345 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_44 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_176 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_175 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_174 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_173 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_344 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_343 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_172 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_344 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_343 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_342 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_341 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_171 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_342 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_341 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_340 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_339 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_170 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_340 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_339 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_338 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_337 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_169 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_338 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_337 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_43 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_172 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_171 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_170 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_169 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_336 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_335 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_168 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_336 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_335 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_334 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_333 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_167 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_334 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_333 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_332 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_331 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_166 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_332 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_331 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_330 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_329 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_165 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_330 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_329 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_42 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_168 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_167 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_166 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_165 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_328 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_327 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_164 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_328 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_327 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_326 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_325 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_163 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_326 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_325 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_324 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_323 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_162 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_324 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_323 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_322 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_321 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_161 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_322 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_321 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_41 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_164 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_163 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_162 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_161 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_11 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_44 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_43 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_42 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_41 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_320 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_319 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_160 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_320 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_319 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_318 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_317 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_159 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_318 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_317 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_316 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_315 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_158 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_316 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_315 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_314 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_313 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_157 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_314 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_313 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_40 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_160 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_159 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_158 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_157 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_312 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_311 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_156 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_312 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_311 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_310 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_309 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_155 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_310 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_309 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_308 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_307 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_154 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_308 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_307 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_306 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_305 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_153 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_306 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_305 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_39 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_156 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_155 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_154 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_153 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_304 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_303 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_152 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_304 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_303 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_302 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_301 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_151 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_302 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_301 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_300 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_299 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_150 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_300 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_299 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_298 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_297 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_149 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_298 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_297 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_38 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_152 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_151 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_150 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_149 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_296 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_295 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_148 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_296 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_295 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_294 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_293 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_147 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_294 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_293 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_292 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_291 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_146 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_292 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_291 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_290 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_289 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_145 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_290 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_289 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_37 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_148 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_147 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_146 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_145 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_10 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  bit2_40 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_39 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_38 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_37 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  CANR2X1 U5 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U10 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_288 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_287 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_144 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_288 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_287 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_286 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_285 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_143 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_286 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_285 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_284 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_283 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_142 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_284 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_283 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_282 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_281 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_141 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_282 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_281 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_36 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_144 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_143 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_142 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_141 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_280 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_279 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_140 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_280 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_279 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_278 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_277 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_139 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_278 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_277 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_276 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_275 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_138 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_276 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_275 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_274 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_273 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_137 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_274 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_273 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_35 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_140 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_139 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_138 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_137 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_272 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_271 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_136 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_272 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_271 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_270 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_269 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_135 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_270 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_269 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_268 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_267 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_134 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_268 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_267 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_266 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_265 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_133 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_266 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_265 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_34 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_136 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_135 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_134 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_133 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_264 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_263 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_132 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_264 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_263 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_262 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_261 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_131 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_262 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_261 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_260 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_259 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_130 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_260 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_259 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_258 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_257 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_129 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_258 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_257 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_33 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_132 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_131 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_130 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_129 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_9 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_36 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_35 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_34 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_33 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_3 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U6 ( .A(s84[3]), .B(n1), .C(s83[3]), .D(n2), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n1), .C(s83[2]), .D(n2), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n1), .C(s83[1]), .D(n2), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n1), .C(s83[0]), .D(n2), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n3), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n3), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n3), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n3), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n1), .C(c_out810), .D(n2), .Z(c_out8) );
  bit4_12 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_11 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_10 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_9 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVDX1 U3 ( .A(n5), .Z0(n1), .Z1(n2) );
  CANR2X1 U4 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n3), .Z(n5) );
  CIVX2 U5 ( .A(c_in8), .Z(n3) );
endmodule


module Add_half_256 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_255 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_128 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_256 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_255 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_254 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_253 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_127 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_254 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_253 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_252 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_251 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_126 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_252 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_251 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_250 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_249 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_125 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_250 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_249 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_32 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_128 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_127 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_126 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_125 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CAOR2XL U4 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U5 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_248 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_247 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_124 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_248 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_247 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_246 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_245 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_123 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_246 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_245 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_244 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_243 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_122 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_244 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_243 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_242 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_241 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_121 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_242 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_241 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_31 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_124 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_123 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_122 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_121 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_240 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_239 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_120 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_240 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_239 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_238 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_237 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_119 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_238 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_237 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_236 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_235 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_118 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_236 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_235 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_234 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_233 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_117 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_234 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_233 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_30 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_120 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_119 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_118 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_117 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_232 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_231 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_116 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_232 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_231 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_230 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_229 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_115 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_230 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_229 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_228 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_227 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_114 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_228 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_227 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_226 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_225 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_113 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_226 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_225 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_29 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_116 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_115 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_114 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_113 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_8 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_32 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_31 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_30 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_29 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_224 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_223 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_112 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_224 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_223 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_222 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_221 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_111 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_222 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_221 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_220 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_219 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_110 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_220 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_219 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_218 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_217 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_109 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_218 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_217 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_28 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_112 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_111 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_110 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_109 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_216 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_215 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_108 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_216 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_215 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_214 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_213 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_107 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_214 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_213 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_212 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_211 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_106 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_212 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_211 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_210 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_209 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_105 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_210 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_209 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_27 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_108 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_107 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_106 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_105 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_208 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_207 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_104 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_208 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_207 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_206 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_205 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_103 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_206 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_205 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_204 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_203 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_102 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_204 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_203 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_202 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_201 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_101 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_202 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_201 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_26 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_104 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_103 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_102 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_101 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_200 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_199 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_100 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_200 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_199 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_198 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_197 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_99 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_198 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_197 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_196 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_195 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_98 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_196 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_195 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_194 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_193 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_97 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_194 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_193 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_25 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_100 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_99 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_98 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_97 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_7 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_28 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_27 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_26 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_25 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_192 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_191 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_96 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_192 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_191 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_190 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_189 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_95 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_190 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_189 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_188 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_187 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_94 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_188 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_187 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_186 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_185 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_93 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_186 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_185 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_24 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_96 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_95 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_94 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_93 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_184 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_183 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_92 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_184 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_183 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_182 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_181 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_91 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_182 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_181 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_180 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_179 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_90 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_180 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_179 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_178 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_177 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_89 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_178 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_177 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_23 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_92 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_91 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_90 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_89 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_176 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_175 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_88 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_176 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_175 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_174 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_173 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_87 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_174 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_173 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_172 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_171 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_86 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_172 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_171 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_170 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_169 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_85 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_170 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_169 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_22 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_88 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_87 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_86 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_85 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_168 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_167 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_84 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_168 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_167 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_166 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_165 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_83 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_166 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_165 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_164 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_163 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_82 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_164 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_163 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_162 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_161 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_81 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_162 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_161 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_21 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_84 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_83 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_82 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_81 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_6 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_24 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_23 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_22 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_21 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_160 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_159 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_80 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_160 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_159 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_158 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_157 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_79 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_158 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_157 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_156 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_155 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_78 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_156 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_155 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_154 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_153 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_77 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_154 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_153 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_20 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_80 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_79 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_78 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_77 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_152 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_151 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_76 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_152 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_151 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_150 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_149 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_75 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_150 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_149 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_148 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_147 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_74 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_148 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_147 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_146 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_145 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_73 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_146 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_145 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_19 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_76 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_75 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_74 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_73 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_144 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_143 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_72 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_144 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_143 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_142 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_141 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_71 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_142 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_141 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_140 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_139 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_70 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_140 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_139 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_138 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_137 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_69 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_138 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_137 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_18 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_72 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_71 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_70 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_69 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_136 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_135 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_68 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_136 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_135 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_134 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_133 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_67 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_134 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_133 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_132 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_131 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_66 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_132 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_131 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_130 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_129 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_65 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_130 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_129 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_17 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_68 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_67 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_66 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_65 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_5 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_20 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_19 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_18 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_17 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_2 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U6 ( .A(s84[3]), .B(n1), .C(s83[3]), .D(n3), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n1), .C(s83[2]), .D(n3), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n1), .C(s83[1]), .D(n3), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n1), .C(s83[0]), .D(n3), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n2), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n2), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n2), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n2), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n1), .C(c_out810), .D(n3), .Z(c_out8) );
  bit4_8 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_7 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_6 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_5 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CANR2X1 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in8), .Z(n2) );
endmodule


module Add_half_128 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_127 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_64 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_128 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_127 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_126 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_125 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_63 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_126 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_125 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_124 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_123 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_62 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_124 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_123 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_122 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_121 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_61 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_122 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_121 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_16 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_64 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_63 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_62 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_61 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_120 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_119 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_60 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_120 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_119 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_118 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_117 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_59 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_118 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_117 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_116 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_115 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_58 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_116 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_115 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_114 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_113 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_57 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_114 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_113 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_15 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_60 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_59 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_58 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_57 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_112 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_111 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_56 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_112 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_111 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_110 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_109 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_55 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_110 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_109 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_108 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_107 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_54 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_108 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_107 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_106 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_105 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_53 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_106 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_105 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_14 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_56 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_55 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_54 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_53 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_104 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_103 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_52 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_104 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_103 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_102 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_101 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_51 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_102 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_101 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_100 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_99 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_50 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_100 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_99 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_98 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_97 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_49 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_98 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_97 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_13 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_52 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_51 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_50 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_49 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_4 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_16 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_15 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_14 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_13 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_96 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_95 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_48 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_96 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_95 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_94 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_93 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_47 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_94 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_93 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_92 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_91 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_46 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_92 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_91 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_90 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_89 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_45 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_90 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_89 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_12 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_48 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_47 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_46 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_45 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_88 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_87 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_44 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_88 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_87 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_86 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_85 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_43 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_86 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_85 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_84 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_83 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_42 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_84 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_83 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_82 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_81 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_41 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_82 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_81 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_11 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_44 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_43 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_42 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_41 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CIVX1 U3 ( .A(n3), .Z(n1) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_80 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_79 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_40 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_80 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_79 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_78 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_77 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_39 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_78 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_77 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_76 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_75 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_38 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_76 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_75 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_74 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_73 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_37 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_74 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_73 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_10 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_40 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_39 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_38 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_37 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_72 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_71 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_36 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_72 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_71 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_70 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_69 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_35 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_70 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_69 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_68 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_67 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_34 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_68 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_67 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_66 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_65 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_33 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_66 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_65 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_9 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_36 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_35 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_34 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_33 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_3 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_12 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_11 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_10 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_9 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_64 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_63 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_32 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_64 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_63 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_62 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_61 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_31 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_62 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_61 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_60 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_59 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_30 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_60 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_59 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_58 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_57 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_29 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_58 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_57 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_8 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_32 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_31 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_30 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_29 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_56 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_55 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_28 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_56 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_55 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_54 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_53 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_27 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_54 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_53 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_52 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_51 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_26 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_52 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_51 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_50 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_49 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_25 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_50 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_49 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_7 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_28 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_27 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_26 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_25 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_48 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_47 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_24 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_48 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_47 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_46 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_45 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_23 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_46 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_45 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_44 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_43 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_22 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_44 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_43 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_42 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_41 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_21 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_42 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_41 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_6 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_24 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_23 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_22 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_21 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_40 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_39 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_20 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_40 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_39 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_38 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_37 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_19 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_38 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_37 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_36 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_35 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_18 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_36 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_35 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_34 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_33 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_17 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_34 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_33 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_5 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_20 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_19 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_18 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_17 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_2 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_8 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_7 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_6 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_5 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_32 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_31 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_16 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_32 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_31 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_30 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_29 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_15 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_30 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_29 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_28 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_27 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_14 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_28 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_27 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_26 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_25 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_13 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_26 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_25 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_4 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_16 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_15 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_14 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_13 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_24 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_23 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_12 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_24 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_23 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_22 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_21 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_11 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_22 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_21 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_20 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_19 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_10 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_20 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_19 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_18 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_17 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_9 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_18 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_17 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_3 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_12 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_11 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_10 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_9 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1)
         );
  CAOR2XL U3 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CANR2X1 U4 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U5 ( .A(n3), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_16 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_15 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_8 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_16 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_15 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_14 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_13 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_7 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_14 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_13 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_12 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_11 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_6 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_12 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_11 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_10 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_9 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_5 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_10 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_9 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_2 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_8 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0)
         );
  Add_full_7 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1)
         );
  Add_full_6 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0)
         );
  Add_full_5 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1)
         );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_8 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_4 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_8 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_6 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_6 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_4 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_4 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module Add_half_2 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
  Add_half_2 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
endmodule


module bit2_1 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  CAOR2X1 U6 ( .A(s4), .B(n1), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n1), .C(c_out10), .D(n3), .Z(c_out2) );
  Add_full_4 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0)
         );
  Add_full_3 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1)
         );
  Add_full_2 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0)
         );
  Add_full_1 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1)
         );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n2) );
endmodule


module bit4_1 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  CAOR2X1 U6 ( .A(s44[1]), .B(n1), .C(s43[1]), .D(n3), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n1), .C(s43[0]), .D(n3), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n1), .C(c_out410), .D(n3), .Z(c_out4) );
  bit2_4 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_3 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_2 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_1 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in4), .Z(n2) );
endmodule


module bit8_1 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  CAOR2X1 U6 ( .A(s84[3]), .B(n1), .C(s83[3]), .D(n3), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n1), .C(s83[2]), .D(n3), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n1), .C(s83[1]), .D(n3), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n1), .C(s83[0]), .D(n3), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n2), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n2), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n2), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n2), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n1), .C(c_out810), .D(n3), .Z(c_out8) );
  bit4_4 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_3 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_2 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_1 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CANR2X1 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CIVX2 U5 ( .A(c_in8), .Z(n2) );
endmodule


module bit16_1 ( sum16, c_out16, a16, b16, c_in16 );
  output [15:0] sum16;
  input [15:0] a16;
  input [15:0] b16;
  input c_in16;
  output c_out16;
  wire   c_out1600, c_out1601, c_out1610, c_out1611, n1, n2, n3, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36;
  wire   [7:0] s161;
  wire   [7:0] s162;
  wire   [7:0] s163;
  wire   [7:0] s164;

  CAOR2X1 U6 ( .A(s164[1]), .B(n34), .C(s163[1]), .D(n36), .Z(sum16[9]) );
  CAOR2X1 U7 ( .A(s164[0]), .B(n34), .C(s163[0]), .D(n36), .Z(sum16[8]) );
  CAOR2X1 U8 ( .A(s162[7]), .B(c_in16), .C(s161[7]), .D(n35), .Z(sum16[7]) );
  CAOR2X1 U9 ( .A(s162[6]), .B(c_in16), .C(s161[6]), .D(n35), .Z(sum16[6]) );
  CAOR2X1 U10 ( .A(s162[5]), .B(c_in16), .C(s161[5]), .D(n35), .Z(sum16[5]) );
  CAOR2X1 U11 ( .A(s162[4]), .B(c_in16), .C(s161[4]), .D(n35), .Z(sum16[4]) );
  CAOR2X1 U12 ( .A(s162[3]), .B(c_in16), .C(s161[3]), .D(n35), .Z(sum16[3]) );
  CAOR2X1 U13 ( .A(s162[2]), .B(c_in16), .C(s161[2]), .D(n35), .Z(sum16[2]) );
  CAOR2X1 U14 ( .A(s162[1]), .B(c_in16), .C(s161[1]), .D(n35), .Z(sum16[1]) );
  CAOR2X1 U15 ( .A(s164[7]), .B(n34), .C(s163[7]), .D(n36), .Z(sum16[15]) );
  CAOR2X1 U16 ( .A(s164[6]), .B(n34), .C(s163[6]), .D(n36), .Z(sum16[14]) );
  CAOR2X1 U17 ( .A(s164[5]), .B(n34), .C(s163[5]), .D(n36), .Z(sum16[13]) );
  CAOR2X1 U18 ( .A(s164[4]), .B(n34), .C(s163[4]), .D(n36), .Z(sum16[12]) );
  CAOR2X1 U19 ( .A(s164[3]), .B(n34), .C(s163[3]), .D(n36), .Z(sum16[11]) );
  CAOR2X1 U20 ( .A(s164[2]), .B(n34), .C(s163[2]), .D(n36), .Z(sum16[10]) );
  CAOR2X1 U21 ( .A(s162[0]), .B(c_in16), .C(s161[0]), .D(n35), .Z(sum16[0]) );
  bit8_4 A161 ( .sum8(s161), .c_out8(c_out1600), .a8({n25, n24, n23, n22, n21, 
        n20, n19, n1}), .b8({n10, n9, n8, n7, n2, n6, n5, n3}), .c_in8(1'b0)
         );
  bit8_3 A162 ( .sum8(s162), .c_out8(c_out1601), .a8({n25, n24, n23, n22, n21, 
        n20, n19, n1}), .b8({n10, n9, n8, n7, n2, n6, n5, n3}), .c_in8(1'b1)
         );
  bit8_2 A163 ( .sum8(s163), .c_out8(c_out1610), .a8({n33, n32, n31, n30, n29, 
        n28, n27, n26}), .b8({n18, n17, n16, n15, n14, n13, n12, n11}), 
        .c_in8(1'b0) );
  bit8_1 A164 ( .sum8(s164), .c_out8(c_out1611), .a8({n33, n32, n31, n30, n29, 
        n28, n27, n26}), .b8({n18, n17, n16, n15, n14, n13, n12, n11}), 
        .c_in8(1'b1) );
  CNIVX3 U3 ( .A(b16[0]), .Z(n3) );
  CNIVX2 U4 ( .A(a16[4]), .Z(n22) );
  CNIVX2 U5 ( .A(b16[2]), .Z(n6) );
  CNIVX2 U22 ( .A(b16[4]), .Z(n7) );
  CNIVX1 U23 ( .A(a16[8]), .Z(n26) );
  CNIVX3 U24 ( .A(a16[0]), .Z(n1) );
  CIVX4 U25 ( .A(n36), .Z(n34) );
  CANR2X4 U26 ( .A(c_out1601), .B(c_in16), .C(c_out1600), .D(n35), .Z(n36) );
  CNIVX2 U27 ( .A(b16[1]), .Z(n5) );
  CNIVX1 U28 ( .A(b16[8]), .Z(n11) );
  CNIVX1 U29 ( .A(b16[5]), .Z(n8) );
  CNIVX1 U30 ( .A(b16[6]), .Z(n9) );
  CNIVX1 U31 ( .A(b16[3]), .Z(n2) );
  CNIVX1 U32 ( .A(b16[12]), .Z(n15) );
  CAOR2XL U33 ( .A(c_out1611), .B(n34), .C(c_out1610), .D(n36), .Z(c_out16) );
  CNIVX1 U34 ( .A(a16[12]), .Z(n30) );
  CNIVX1 U35 ( .A(a16[3]), .Z(n21) );
  CNIVX1 U36 ( .A(a16[1]), .Z(n19) );
  CNIVX1 U37 ( .A(a16[2]), .Z(n20) );
  CNIVX1 U38 ( .A(b16[13]), .Z(n16) );
  CNIVX1 U39 ( .A(b16[7]), .Z(n10) );
  CNIVX1 U40 ( .A(b16[14]), .Z(n17) );
  CNIVX1 U41 ( .A(b16[11]), .Z(n14) );
  CNIVX1 U42 ( .A(b16[10]), .Z(n13) );
  CNIVX1 U43 ( .A(b16[9]), .Z(n12) );
  CNIVX1 U44 ( .A(b16[15]), .Z(n18) );
  CNIVX1 U45 ( .A(a16[7]), .Z(n25) );
  CNIVX1 U46 ( .A(a16[11]), .Z(n29) );
  CNIVX1 U47 ( .A(a16[13]), .Z(n31) );
  CNIVX1 U48 ( .A(a16[14]), .Z(n32) );
  CNIVX1 U49 ( .A(a16[15]), .Z(n33) );
  CNIVX1 U50 ( .A(a16[5]), .Z(n23) );
  CNIVX1 U51 ( .A(a16[6]), .Z(n24) );
  CNIVX1 U52 ( .A(a16[9]), .Z(n27) );
  CNIVX1 U53 ( .A(a16[10]), .Z(n28) );
  CIVX2 U54 ( .A(c_in16), .Z(n35) );
endmodule


module bit32 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   c_out3200, c_out3201, c_out3210, c_out3211, n4, n1, n2, n3, n5, n6;
  wire   [15:0] s321;
  wire   [15:0] s322;
  wire   [15:0] s323;
  wire   [15:0] s324;

  CAOR2X1 U6 ( .A(s322[9]), .B(c_in32), .C(s321[9]), .D(n6), .Z(sum32[9]) );
  CAOR2X1 U7 ( .A(s322[8]), .B(c_in32), .C(s321[8]), .D(n6), .Z(sum32[8]) );
  CAOR2X1 U8 ( .A(s322[7]), .B(c_in32), .C(s321[7]), .D(n6), .Z(sum32[7]) );
  CAOR2X1 U9 ( .A(s322[6]), .B(c_in32), .C(s321[6]), .D(n6), .Z(sum32[6]) );
  CAOR2X1 U10 ( .A(s322[5]), .B(c_in32), .C(s321[5]), .D(n6), .Z(sum32[5]) );
  CAOR2X1 U11 ( .A(s322[4]), .B(c_in32), .C(s321[4]), .D(n6), .Z(sum32[4]) );
  CAOR2X1 U12 ( .A(s322[3]), .B(c_in32), .C(s321[3]), .D(n6), .Z(sum32[3]) );
  CAOR2X1 U13 ( .A(s324[15]), .B(n5), .C(s323[15]), .D(n3), .Z(sum32[31]) );
  CAOR2X1 U14 ( .A(s324[14]), .B(n5), .C(s323[14]), .D(n3), .Z(sum32[30]) );
  CAOR2X1 U15 ( .A(s322[2]), .B(c_in32), .C(s321[2]), .D(n6), .Z(sum32[2]) );
  CAOR2X1 U16 ( .A(s324[13]), .B(n5), .C(s323[13]), .D(n3), .Z(sum32[29]) );
  CAOR2X1 U17 ( .A(s324[12]), .B(n5), .C(s323[12]), .D(n3), .Z(sum32[28]) );
  CAOR2X1 U18 ( .A(s324[11]), .B(n5), .C(s323[11]), .D(n3), .Z(sum32[27]) );
  CAOR2X1 U19 ( .A(s324[10]), .B(n5), .C(s323[10]), .D(n3), .Z(sum32[26]) );
  CAOR2X1 U22 ( .A(s324[7]), .B(n5), .C(s323[7]), .D(n3), .Z(sum32[23]) );
  CAOR2X1 U23 ( .A(s324[6]), .B(n5), .C(s323[6]), .D(n3), .Z(sum32[22]) );
  CAOR2X1 U24 ( .A(s324[5]), .B(n5), .C(s323[5]), .D(n3), .Z(sum32[21]) );
  CAOR2X1 U25 ( .A(s324[4]), .B(n5), .C(s323[4]), .D(n3), .Z(sum32[20]) );
  CAOR2X1 U26 ( .A(s322[1]), .B(c_in32), .C(s321[1]), .D(n6), .Z(sum32[1]) );
  CAOR2X1 U31 ( .A(s322[15]), .B(c_in32), .C(s321[15]), .D(n6), .Z(sum32[15])
         );
  CAOR2X1 U32 ( .A(s322[14]), .B(c_in32), .C(s321[14]), .D(n6), .Z(sum32[14])
         );
  CAOR2X1 U33 ( .A(s322[13]), .B(c_in32), .C(s321[13]), .D(n6), .Z(sum32[13])
         );
  CAOR2X1 U34 ( .A(s322[12]), .B(c_in32), .C(s321[12]), .D(n6), .Z(sum32[12])
         );
  CAOR2X1 U35 ( .A(s322[11]), .B(c_in32), .C(s321[11]), .D(n6), .Z(sum32[11])
         );
  CAOR2X1 U36 ( .A(s322[10]), .B(c_in32), .C(s321[10]), .D(n6), .Z(sum32[10])
         );
  CAOR2X1 U37 ( .A(s322[0]), .B(c_in32), .C(s321[0]), .D(n6), .Z(sum32[0]) );
  bit16_0 A321 ( .sum16(s321), .c_out16(c_out3200), .a16(a32[15:0]), .b16(
        b32[15:0]), .c_in16(1'b0) );
  bit16_3 A322 ( .sum16(s322), .c_out16(c_out3201), .a16(a32[15:0]), .b16(
        b32[15:0]), .c_in16(1'b1) );
  bit16_2 A323 ( .sum16(s323), .c_out16(c_out3210), .a16(a32[31:16]), .b16(
        b32[31:16]), .c_in16(1'b0) );
  bit16_1 A324 ( .sum16(s324), .c_out16(c_out3211), .a16(a32[31:16]), .b16(
        b32[31:16]), .c_in16(1'b1) );
  CND2X1 U3 ( .A(c_out3201), .B(c_in32), .Z(n1) );
  CND2X1 U4 ( .A(c_out3200), .B(n6), .Z(n2) );
  CIVDX3 U5 ( .A(n4), .Z0(n5), .Z1(n3) );
  CAN2X2 U20 ( .A(n1), .B(n2), .Z(n4) );
  CAOR2XL U21 ( .A(s324[9]), .B(n5), .C(s323[9]), .D(n3), .Z(sum32[25]) );
  CAOR2XL U27 ( .A(s324[8]), .B(n5), .C(s323[8]), .D(n3), .Z(sum32[24]) );
  CAOR2XL U28 ( .A(s324[1]), .B(n5), .C(s323[1]), .D(n3), .Z(sum32[17]) );
  CAOR2XL U29 ( .A(s324[2]), .B(n5), .C(s323[2]), .D(n3), .Z(sum32[18]) );
  CAOR2XL U30 ( .A(s324[3]), .B(n5), .C(s323[3]), .D(n3), .Z(sum32[19]) );
  CAOR2XL U38 ( .A(s324[0]), .B(n5), .C(s323[0]), .D(n3), .Z(sum32[16]) );
  CAOR2XL U39 ( .A(n5), .B(c_out3211), .C(c_out3210), .D(n3), .Z(c_out32) );
  CIVX2 U40 ( .A(c_in32), .Z(n6) );
endmodule


module seq_adder_DW01_dec_1 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n5, n6, n7, n8, n9, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n34, n36, n37, n38, n40, n41, n43, n44,
         n45, n47, n50, n51, n53, n54, n57, n60, n61, n64, n68, n69, n71, n72,
         n73, n75, n77, n79, n80, n81, n82, n84, n86, n88, n90, n91, n92, n94,
         n96, n98, n99, n100, n103, n106, n107, n108, n109, n112, n115, n116,
         n119, n123, n124, n125, n128, n131, n132, n135, n205;
  assign n1 = A[24];
  assign n5 = A[20];
  assign n6 = A[19];
  assign n7 = A[18];
  assign n8 = A[17];
  assign n9 = A[16];
  assign n16 = A[9];
  assign n17 = A[8];
  assign n18 = A[7];
  assign n19 = A[6];
  assign n20 = A[5];
  assign n21 = A[4];
  assign n22 = A[3];
  assign n23 = A[2];
  assign n24 = A[1];
  assign n38 = A[23];
  assign n41 = A[22];
  assign n45 = A[21];
  assign n73 = A[15];
  assign n77 = A[14];
  assign n82 = A[13];
  assign n86 = A[12];
  assign n92 = A[11];
  assign n96 = A[10];
  assign n135 = A[0];

  COR2X1 U3 ( .A(A[30]), .B(n26), .Z(n25) );
  COR2X1 U5 ( .A(A[29]), .B(n27), .Z(n26) );
  COR2X1 U7 ( .A(A[28]), .B(n28), .Z(n27) );
  COR2X1 U9 ( .A(A[27]), .B(n29), .Z(n28) );
  COR2X1 U11 ( .A(A[26]), .B(n30), .Z(n29) );
  COR2X1 U13 ( .A(A[25]), .B(n205), .Z(n30) );
  COR2X1 U171 ( .A(n69), .B(n53), .Z(n51) );
  COR4X1 U172 ( .A(n124), .B(n108), .C(n71), .D(n90), .Z(n69) );
  COR2X1 U173 ( .A(n106), .B(n90), .Z(n88) );
  COR2X1 U174 ( .A(n69), .B(n9), .Z(n64) );
  COR3X2 U175 ( .A(n106), .B(n90), .C(n86), .Z(n84) );
  COR3X2 U176 ( .A(n69), .B(n53), .C(n36), .Z(n34) );
  COR2X1 U177 ( .A(n124), .B(n21), .Z(n119) );
  COR3X2 U178 ( .A(n88), .B(n80), .C(n77), .Z(n75) );
  COR3X2 U179 ( .A(n106), .B(n99), .C(n96), .Z(n94) );
  COR4X1 U180 ( .A(n69), .B(n53), .C(n36), .D(n1), .Z(n205) );
  CNR2X1 U181 ( .A(n88), .B(n80), .Z(n79) );
  CNR2X1 U182 ( .A(n106), .B(n99), .Z(n98) );
  CND2X1 U183 ( .A(n50), .B(n44), .Z(n43) );
  CND2X1 U184 ( .A(n68), .B(n61), .Z(n60) );
  CND2X1 U185 ( .A(n123), .B(n116), .Z(n115) );
  CNR2X1 U186 ( .A(n20), .B(n21), .Z(n116) );
  CNR2X1 U187 ( .A(n5), .B(n45), .Z(n44) );
  CNR2X1 U188 ( .A(n9), .B(n8), .Z(n61) );
  CND2X1 U189 ( .A(n44), .B(n37), .Z(n36) );
  CNR2X1 U190 ( .A(n41), .B(n38), .Z(n37) );
  CNR2X1 U191 ( .A(n135), .B(n24), .Z(n132) );
  CNR2X1 U192 ( .A(n17), .B(n16), .Z(n100) );
  CNR2X1 U193 ( .A(n86), .B(n82), .Z(n81) );
  CNR2X1 U194 ( .A(n124), .B(n108), .Z(n107) );
  CND2X1 U195 ( .A(n116), .B(n109), .Z(n108) );
  CNR2X1 U196 ( .A(n19), .B(n18), .Z(n109) );
  CND2X1 U197 ( .A(n100), .B(n91), .Z(n90) );
  CNR2X1 U198 ( .A(n92), .B(n96), .Z(n91) );
  CND2X1 U199 ( .A(n132), .B(n125), .Z(n124) );
  CNR2X1 U200 ( .A(n23), .B(n22), .Z(n125) );
  CND2X1 U201 ( .A(n61), .B(n54), .Z(n53) );
  CNR2X1 U202 ( .A(n7), .B(n6), .Z(n54) );
  CND2X1 U203 ( .A(n81), .B(n72), .Z(n71) );
  CNR2X1 U204 ( .A(n77), .B(n73), .Z(n72) );
  CENX1 U205 ( .A(A[30]), .B(n26), .Z(SUM[30]) );
  CENX1 U206 ( .A(A[29]), .B(n27), .Z(SUM[29]) );
  CENX1 U207 ( .A(A[28]), .B(n28), .Z(SUM[28]) );
  CENX1 U208 ( .A(A[31]), .B(n25), .Z(SUM[31]) );
  CNR2X1 U209 ( .A(n43), .B(n41), .Z(n40) );
  CNR2X1 U210 ( .A(n51), .B(n5), .Z(n47) );
  CNR2X1 U211 ( .A(n60), .B(n7), .Z(n57) );
  CNR2X1 U212 ( .A(n106), .B(n17), .Z(n103) );
  CNR2X1 U213 ( .A(n115), .B(n19), .Z(n112) );
  CEOX1 U214 ( .A(n21), .B(n123), .Z(SUM[4]) );
  CEOX1 U215 ( .A(n22), .B(n128), .Z(SUM[3]) );
  CENX1 U216 ( .A(n131), .B(n23), .Z(SUM[2]) );
  CENX1 U217 ( .A(n135), .B(n24), .Z(SUM[1]) );
  CENX1 U218 ( .A(n119), .B(n20), .Z(SUM[5]) );
  CENX1 U219 ( .A(A[27]), .B(n29), .Z(SUM[27]) );
  CENX1 U220 ( .A(A[26]), .B(n30), .Z(SUM[26]) );
  CENX1 U221 ( .A(A[25]), .B(n205), .Z(SUM[25]) );
  CENX1 U222 ( .A(n34), .B(n1), .Z(SUM[24]) );
  CEOX1 U223 ( .A(n38), .B(n40), .Z(SUM[23]) );
  CENX1 U224 ( .A(n43), .B(n41), .Z(SUM[22]) );
  CEOX1 U225 ( .A(n45), .B(n47), .Z(SUM[21]) );
  CEOX1 U226 ( .A(n5), .B(n50), .Z(SUM[20]) );
  CEOX1 U227 ( .A(n6), .B(n57), .Z(SUM[19]) );
  CENX1 U228 ( .A(n60), .B(n7), .Z(SUM[18]) );
  CENX1 U229 ( .A(n64), .B(n8), .Z(SUM[17]) );
  CEOX1 U230 ( .A(n9), .B(n68), .Z(SUM[16]) );
  CENX1 U231 ( .A(n75), .B(n73), .Z(SUM[15]) );
  CEOX1 U232 ( .A(n77), .B(n79), .Z(SUM[14]) );
  CENX1 U233 ( .A(n84), .B(n82), .Z(SUM[13]) );
  CENX1 U234 ( .A(n88), .B(n86), .Z(SUM[12]) );
  CENX1 U235 ( .A(n94), .B(n92), .Z(SUM[11]) );
  CEOX1 U236 ( .A(n96), .B(n98), .Z(SUM[10]) );
  CEOX1 U237 ( .A(n16), .B(n103), .Z(SUM[9]) );
  CEOX1 U238 ( .A(n18), .B(n112), .Z(SUM[7]) );
  CNR2X1 U239 ( .A(n131), .B(n23), .Z(n128) );
  CENX1 U240 ( .A(n106), .B(n17), .Z(SUM[8]) );
  CENX1 U241 ( .A(n115), .B(n19), .Z(SUM[6]) );
  CIVX2 U242 ( .A(n100), .Z(n99) );
  CIVX2 U243 ( .A(n81), .Z(n80) );
  CIVX2 U244 ( .A(n69), .Z(n68) );
  CIVX2 U245 ( .A(n51), .Z(n50) );
  CIVX2 U246 ( .A(n132), .Z(n131) );
  CIVX2 U247 ( .A(n124), .Z(n123) );
  CIVX2 U248 ( .A(n107), .Z(n106) );
  CIVX2 U249 ( .A(n135), .Z(SUM[0]) );
endmodule


module seq_adder ( clock, start, valid, mlier, mcand, prodt_end, reset );
  input [31:0] mlier;
  input [31:0] mcand;
  output [64:0] prodt_end;
  input clock, start, reset;
  output valid;
  wire   wcout, add, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N326, N327, n12, n13, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n163,
         n164, n165, n166, n167, n169, n170, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n419,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567;
  wire   [31:0] a;
  wire   [31:0] wsum;
  wire   [1:0] states;
  wire   [31:0] count;
  wire   [31:0] b;
  assign prodt_end[64] = 1'b0;

  CAOR1X1 U306 ( .A(prodt_end[0]), .B(n415), .C(n161), .Z(n315) );
  CAOR2X1 U307 ( .A(n525), .B(a[31]), .C(n531), .D(mcand[31]), .Z(n316) );
  CAOR2X1 U308 ( .A(n525), .B(a[30]), .C(n531), .D(mcand[30]), .Z(n317) );
  CAOR2X1 U309 ( .A(n525), .B(a[29]), .C(n531), .D(mcand[29]), .Z(n318) );
  CAOR2X1 U310 ( .A(n525), .B(a[28]), .C(n531), .D(mcand[28]), .Z(n319) );
  CAOR2X1 U311 ( .A(n525), .B(a[27]), .C(n531), .D(mcand[27]), .Z(n320) );
  CAOR2X1 U312 ( .A(n525), .B(a[26]), .C(n531), .D(mcand[26]), .Z(n321) );
  CAOR2X1 U313 ( .A(n525), .B(a[25]), .C(n531), .D(mcand[25]), .Z(n322) );
  CAOR2X1 U314 ( .A(n525), .B(a[24]), .C(n531), .D(mcand[24]), .Z(n323) );
  CAOR2X1 U315 ( .A(n525), .B(a[23]), .C(n531), .D(mcand[23]), .Z(n324) );
  CAOR2X1 U316 ( .A(n525), .B(a[22]), .C(n531), .D(mcand[22]), .Z(n325) );
  CAOR2X1 U317 ( .A(n525), .B(a[21]), .C(n531), .D(mcand[21]), .Z(n326) );
  CAOR2X1 U318 ( .A(n525), .B(a[20]), .C(n531), .D(mcand[20]), .Z(n327) );
  CAOR2X1 U319 ( .A(n525), .B(a[19]), .C(n531), .D(mcand[19]), .Z(n328) );
  CAOR2X1 U320 ( .A(n525), .B(a[18]), .C(n531), .D(mcand[18]), .Z(n329) );
  CAOR2X1 U321 ( .A(n525), .B(a[17]), .C(n531), .D(mcand[17]), .Z(n330) );
  CAOR2X1 U322 ( .A(n525), .B(a[16]), .C(n531), .D(mcand[16]), .Z(n331) );
  CAOR2X1 U323 ( .A(n525), .B(a[15]), .C(n531), .D(mcand[15]), .Z(n332) );
  CAOR2X1 U324 ( .A(n525), .B(a[14]), .C(n531), .D(mcand[14]), .Z(n333) );
  CAOR2X1 U325 ( .A(n525), .B(a[13]), .C(n531), .D(mcand[13]), .Z(n334) );
  CAOR2X1 U326 ( .A(n525), .B(a[12]), .C(n531), .D(mcand[12]), .Z(n335) );
  CAOR2X1 U327 ( .A(n525), .B(a[11]), .C(n531), .D(mcand[11]), .Z(n336) );
  CAOR2X1 U329 ( .A(n525), .B(a[9]), .C(n531), .D(mcand[9]), .Z(n338) );
  CAOR2X1 U331 ( .A(n525), .B(a[7]), .C(n531), .D(mcand[7]), .Z(n340) );
  CAOR2X1 U334 ( .A(n525), .B(a[4]), .C(n531), .D(mcand[4]), .Z(n343) );
  CAOR2X1 U339 ( .A(n525), .B(b[30]), .C(mlier[30]), .D(n531), .Z(n349) );
  CAOR2X1 U340 ( .A(n525), .B(b[29]), .C(mlier[29]), .D(n531), .Z(n350) );
  CAOR2X1 U341 ( .A(n525), .B(b[28]), .C(mlier[28]), .D(n531), .Z(n351) );
  CAOR2X1 U342 ( .A(n525), .B(b[27]), .C(mlier[27]), .D(n531), .Z(n352) );
  CAOR2X1 U343 ( .A(n525), .B(b[26]), .C(mlier[26]), .D(n531), .Z(n353) );
  CAOR2X1 U344 ( .A(n525), .B(b[25]), .C(mlier[25]), .D(n531), .Z(n354) );
  CAOR2X1 U345 ( .A(n525), .B(b[24]), .C(mlier[24]), .D(n531), .Z(n355) );
  CAOR2X1 U346 ( .A(n525), .B(b[23]), .C(mlier[23]), .D(n531), .Z(n356) );
  CAOR2X1 U347 ( .A(n525), .B(b[22]), .C(mlier[22]), .D(n531), .Z(n357) );
  CAOR2X1 U348 ( .A(n525), .B(b[21]), .C(mlier[21]), .D(n531), .Z(n358) );
  CAOR2X1 U349 ( .A(n525), .B(b[20]), .C(mlier[20]), .D(n531), .Z(n359) );
  CAOR2X1 U350 ( .A(n525), .B(b[19]), .C(mlier[19]), .D(n531), .Z(n360) );
  CAOR2X1 U351 ( .A(n525), .B(b[18]), .C(mlier[18]), .D(n531), .Z(n361) );
  CAOR2X1 U352 ( .A(n525), .B(b[17]), .C(mlier[17]), .D(n531), .Z(n362) );
  CAOR2X1 U353 ( .A(n525), .B(b[16]), .C(mlier[16]), .D(n531), .Z(n363) );
  CAOR2X1 U354 ( .A(n525), .B(b[15]), .C(mlier[15]), .D(n531), .Z(n364) );
  CAOR2X1 U355 ( .A(n525), .B(b[14]), .C(mlier[14]), .D(n531), .Z(n365) );
  CAOR2X1 U356 ( .A(n525), .B(b[13]), .C(mlier[13]), .D(n531), .Z(n366) );
  CAOR2X1 U357 ( .A(n525), .B(b[12]), .C(mlier[12]), .D(n531), .Z(n367) );
  CAOR2X1 U358 ( .A(n525), .B(b[11]), .C(mlier[11]), .D(n531), .Z(n368) );
  CAOR2X1 U359 ( .A(n525), .B(b[10]), .C(mlier[10]), .D(n531), .Z(n369) );
  CAOR2X1 U360 ( .A(n525), .B(b[9]), .C(mlier[9]), .D(n531), .Z(n370) );
  CAOR2X1 U361 ( .A(n525), .B(b[8]), .C(mlier[8]), .D(n531), .Z(n371) );
  CAOR2X1 U362 ( .A(n525), .B(b[7]), .C(mlier[7]), .D(n531), .Z(n372) );
  CAOR2X1 U363 ( .A(n525), .B(b[6]), .C(mlier[6]), .D(n531), .Z(n373) );
  CAOR2X1 U364 ( .A(n525), .B(b[5]), .C(mlier[5]), .D(n531), .Z(n374) );
  CAOR2X1 U365 ( .A(n525), .B(b[4]), .C(mlier[4]), .D(n531), .Z(n375) );
  CAOR2X1 U366 ( .A(n525), .B(b[3]), .C(mlier[3]), .D(n531), .Z(n376) );
  CAOR2X1 U367 ( .A(n525), .B(b[2]), .C(mlier[2]), .D(n531), .Z(n377) );
  CAOR2X1 U368 ( .A(n525), .B(b[1]), .C(n531), .D(mlier[1]), .Z(n378) );
  CAOR2X1 U400 ( .A(n527), .B(n167), .C(n426), .D(n535), .Z(N327) );
  CNR8X1 U401 ( .A(count[31]), .B(count[3]), .C(count[4]), .D(count[5]), .E(
        count[6]), .F(count[7]), .G(count[8]), .H(count[9]), .Z(n252) );
  CNR8X1 U402 ( .A(count[24]), .B(count[25]), .C(count[26]), .D(count[27]), 
        .E(count[28]), .F(count[29]), .G(count[2]), .H(count[30]), .Z(n251) );
  CNR8X1 U403 ( .A(count[17]), .B(count[18]), .C(count[19]), .D(count[1]), .E(
        count[20]), .F(count[21]), .G(count[22]), .H(count[23]), .Z(n250) );
  CNR8X1 U404 ( .A(n519), .B(count[10]), .C(count[11]), .D(count[12]), .E(
        count[13]), .F(count[14]), .G(count[15]), .H(count[16]), .Z(n249) );
  bit32 Ad32 ( .a32(prodt_end[63:32]), .b32(a), .sum32(wsum), .c_out32(wcout), 
        .c_in32(1'b0) );
  seq_adder_DW01_dec_1 sub_72 ( .A(count), .SUM({N86, N85, N84, N83, N82, N81, 
        N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, 
        N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55}) );
  CFD1QX4 \prodt_end_reg[32]  ( .D(n284), .CP(clock), .Q(prodt_end[32]) );
  CFD1QXL \prodt_end_reg[31]  ( .D(n285), .CP(clock), .Q(prodt_end[31]) );
  CFD1QX1 \a_reg[24]  ( .D(n323), .CP(clock), .Q(a[24]) );
  CFD1QX4 \a_reg[0]  ( .D(n347), .CP(clock), .Q(a[0]) );
  CFD1QXL \prodt_end_reg[0]  ( .D(n315), .CP(clock), .Q(prodt_end[0]) );
  CFD1QXL \prodt_end_reg[1]  ( .D(n413), .CP(clock), .Q(prodt_end[1]) );
  CFD1QXL \prodt_end_reg[30]  ( .D(n286), .CP(clock), .Q(prodt_end[30]) );
  CFD1QXL \prodt_end_reg[29]  ( .D(n287), .CP(clock), .Q(prodt_end[29]) );
  CFD1QXL \prodt_end_reg[28]  ( .D(n288), .CP(clock), .Q(prodt_end[28]) );
  CFD1QXL \prodt_end_reg[27]  ( .D(n289), .CP(clock), .Q(prodt_end[27]) );
  CFD1QXL \prodt_end_reg[26]  ( .D(n290), .CP(clock), .Q(prodt_end[26]) );
  CFD1QXL \prodt_end_reg[25]  ( .D(n291), .CP(clock), .Q(prodt_end[25]) );
  CFD1QXL \prodt_end_reg[24]  ( .D(n292), .CP(clock), .Q(prodt_end[24]) );
  CFD1QXL \prodt_end_reg[23]  ( .D(n293), .CP(clock), .Q(prodt_end[23]) );
  CFD1QXL \prodt_end_reg[22]  ( .D(n294), .CP(clock), .Q(prodt_end[22]) );
  CFD1QXL \prodt_end_reg[21]  ( .D(n295), .CP(clock), .Q(prodt_end[21]) );
  CFD1QXL \prodt_end_reg[20]  ( .D(n296), .CP(clock), .Q(prodt_end[20]) );
  CFD1QXL \prodt_end_reg[19]  ( .D(n297), .CP(clock), .Q(prodt_end[19]) );
  CFD1QXL \prodt_end_reg[18]  ( .D(n298), .CP(clock), .Q(prodt_end[18]) );
  CFD1QXL \prodt_end_reg[17]  ( .D(n299), .CP(clock), .Q(prodt_end[17]) );
  CFD1QXL \prodt_end_reg[16]  ( .D(n300), .CP(clock), .Q(prodt_end[16]) );
  CFD1QXL \prodt_end_reg[15]  ( .D(n301), .CP(clock), .Q(prodt_end[15]) );
  CFD1QXL \prodt_end_reg[14]  ( .D(n302), .CP(clock), .Q(prodt_end[14]) );
  CFD1QXL \prodt_end_reg[13]  ( .D(n303), .CP(clock), .Q(prodt_end[13]) );
  CFD1QXL \prodt_end_reg[12]  ( .D(n304), .CP(clock), .Q(prodt_end[12]) );
  CFD1QXL \prodt_end_reg[11]  ( .D(n305), .CP(clock), .Q(prodt_end[11]) );
  CFD1QXL \prodt_end_reg[10]  ( .D(n306), .CP(clock), .Q(prodt_end[10]) );
  CFD1QXL \prodt_end_reg[9]  ( .D(n307), .CP(clock), .Q(prodt_end[9]) );
  CFD1QXL \prodt_end_reg[8]  ( .D(n308), .CP(clock), .Q(prodt_end[8]) );
  CFD1QXL \prodt_end_reg[7]  ( .D(n309), .CP(clock), .Q(prodt_end[7]) );
  CFD1QXL \prodt_end_reg[6]  ( .D(n310), .CP(clock), .Q(prodt_end[6]) );
  CFD1QXL \prodt_end_reg[5]  ( .D(n311), .CP(clock), .Q(prodt_end[5]) );
  CFD1QXL \prodt_end_reg[4]  ( .D(n312), .CP(clock), .Q(prodt_end[4]) );
  CFD1QXL \prodt_end_reg[3]  ( .D(n313), .CP(clock), .Q(prodt_end[3]) );
  CFD1QXL \prodt_end_reg[2]  ( .D(n314), .CP(clock), .Q(prodt_end[2]) );
  CFD1QXL valid_reg ( .D(n380), .CP(clock), .Q(valid) );
  CFD1QXL \b_reg[30]  ( .D(n349), .CP(clock), .Q(b[30]) );
  CFD1QXL \b_reg[29]  ( .D(n350), .CP(clock), .Q(b[29]) );
  CFD1QXL \b_reg[28]  ( .D(n351), .CP(clock), .Q(b[28]) );
  CFD1QXL \b_reg[25]  ( .D(n354), .CP(clock), .Q(b[25]) );
  CFD1QXL \b_reg[24]  ( .D(n355), .CP(clock), .Q(b[24]) );
  CFD1QXL \b_reg[23]  ( .D(n356), .CP(clock), .Q(b[23]) );
  CFD1QXL \b_reg[22]  ( .D(n357), .CP(clock), .Q(b[22]) );
  CFD1QXL \b_reg[21]  ( .D(n358), .CP(clock), .Q(b[21]) );
  CFD1QXL \b_reg[20]  ( .D(n359), .CP(clock), .Q(b[20]) );
  CFD1QXL \b_reg[19]  ( .D(n360), .CP(clock), .Q(b[19]) );
  CFD1QXL \b_reg[18]  ( .D(n361), .CP(clock), .Q(b[18]) );
  CFD1QXL \b_reg[17]  ( .D(n362), .CP(clock), .Q(b[17]) );
  CFD1QXL \b_reg[16]  ( .D(n363), .CP(clock), .Q(b[16]) );
  CFD1QXL \b_reg[15]  ( .D(n364), .CP(clock), .Q(b[15]) );
  CFD1QXL \b_reg[14]  ( .D(n365), .CP(clock), .Q(b[14]) );
  CFD1QXL \b_reg[13]  ( .D(n366), .CP(clock), .Q(b[13]) );
  CFD1QXL \b_reg[12]  ( .D(n367), .CP(clock), .Q(b[12]) );
  CFD1QXL \b_reg[11]  ( .D(n368), .CP(clock), .Q(b[11]) );
  CFD1QXL \b_reg[10]  ( .D(n369), .CP(clock), .Q(b[10]) );
  CFD1QXL \b_reg[9]  ( .D(n370), .CP(clock), .Q(b[9]) );
  CFD1QXL \b_reg[8]  ( .D(n371), .CP(clock), .Q(b[8]) );
  CFD1QXL \b_reg[7]  ( .D(n372), .CP(clock), .Q(b[7]) );
  CFD1QXL \b_reg[6]  ( .D(n373), .CP(clock), .Q(b[6]) );
  CFD1QXL \b_reg[5]  ( .D(n374), .CP(clock), .Q(b[5]) );
  CFD1QXL \b_reg[4]  ( .D(n375), .CP(clock), .Q(b[4]) );
  CFD1QXL \b_reg[3]  ( .D(n376), .CP(clock), .Q(b[3]) );
  CFD1QXL \b_reg[2]  ( .D(n377), .CP(clock), .Q(b[2]) );
  CFD1QXL \b_reg[1]  ( .D(n378), .CP(clock), .Q(b[1]) );
  CFD1QXL \b_reg[27]  ( .D(n352), .CP(clock), .Q(b[27]) );
  CFD1QXL \b_reg[26]  ( .D(n353), .CP(clock), .Q(b[26]) );
  CFD1QXL \count_reg[31]  ( .D(n381), .CP(clock), .Q(count[31]) );
  CFD1QXL \count_reg[30]  ( .D(n382), .CP(clock), .Q(count[30]) );
  CFD1QXL \count_reg[25]  ( .D(n387), .CP(clock), .Q(count[25]) );
  CFD1QXL \count_reg[26]  ( .D(n386), .CP(clock), .Q(count[26]) );
  CFD1QXL \count_reg[29]  ( .D(n383), .CP(clock), .Q(count[29]) );
  CFD1QXL \count_reg[27]  ( .D(n385), .CP(clock), .Q(count[27]) );
  CFD1QXL \count_reg[28]  ( .D(n384), .CP(clock), .Q(count[28]) );
  CFD1XL \b_reg[31]  ( .D(n348), .CP(clock), .QN(n12) );
  CFD1XL \b_reg[0]  ( .D(n379), .CP(clock), .QN(n13) );
  CFD1QXL add_reg ( .D(n414), .CP(clock), .Q(add) );
  CFD1QXL \states_reg[1]  ( .D(N327), .CP(clock), .Q(states[1]) );
  CFD1QXL \states_reg[0]  ( .D(N326), .CP(clock), .Q(states[0]) );
  CFD1XL \count_reg[5]  ( .D(n407), .CP(clock), .Q(count[5]) );
  CFD1QXL \count_reg[24]  ( .D(n388), .CP(clock), .Q(count[24]) );
  CFD1QXL \count_reg[11]  ( .D(n401), .CP(clock), .Q(count[11]) );
  CFD1QXL \count_reg[17]  ( .D(n395), .CP(clock), .Q(count[17]) );
  CFD1QXL \count_reg[15]  ( .D(n397), .CP(clock), .Q(count[15]) );
  CFD1QXL \count_reg[13]  ( .D(n399), .CP(clock), .Q(count[13]) );
  CFD1QXL \count_reg[9]  ( .D(n403), .CP(clock), .Q(count[9]) );
  CFD1QXL \count_reg[23]  ( .D(n389), .CP(clock), .Q(count[23]) );
  CFD1QXL \count_reg[19]  ( .D(n393), .CP(clock), .Q(count[19]) );
  CFD1QXL \count_reg[7]  ( .D(n405), .CP(clock), .Q(count[7]) );
  CFD1QXL \count_reg[21]  ( .D(n391), .CP(clock), .Q(count[21]) );
  CFD1QXL \count_reg[1]  ( .D(n411), .CP(clock), .Q(count[1]) );
  CFD1QXL \count_reg[3]  ( .D(n409), .CP(clock), .Q(count[3]) );
  CFD1QXL \count_reg[12]  ( .D(n400), .CP(clock), .Q(count[12]) );
  CFD1QXL \count_reg[16]  ( .D(n396), .CP(clock), .Q(count[16]) );
  CFD1QXL \count_reg[14]  ( .D(n398), .CP(clock), .Q(count[14]) );
  CFD1QXL \count_reg[18]  ( .D(n394), .CP(clock), .Q(count[18]) );
  CFD1QXL \count_reg[22]  ( .D(n390), .CP(clock), .Q(count[22]) );
  CFD1QXL \count_reg[10]  ( .D(n402), .CP(clock), .Q(count[10]) );
  CFD1QXL \count_reg[20]  ( .D(n392), .CP(clock), .Q(count[20]) );
  CFD1QXL \count_reg[2]  ( .D(n410), .CP(clock), .Q(count[2]) );
  CFD1QXL \count_reg[4]  ( .D(n408), .CP(clock), .Q(count[4]) );
  CFD1QXL \count_reg[8]  ( .D(n404), .CP(clock), .Q(count[8]) );
  CFD1QXL \count_reg[6]  ( .D(n406), .CP(clock), .Q(count[6]) );
  CFD1QXL \prodt_end_reg[63]  ( .D(n253), .CP(clock), .Q(prodt_end[63]) );
  CFD1QXL \prodt_end_reg[62]  ( .D(n254), .CP(clock), .Q(prodt_end[62]) );
  CFD1QXL \prodt_end_reg[61]  ( .D(n255), .CP(clock), .Q(prodt_end[61]) );
  CFD1QXL \prodt_end_reg[58]  ( .D(n258), .CP(clock), .Q(prodt_end[58]) );
  CFD1QXL \prodt_end_reg[57]  ( .D(n259), .CP(clock), .Q(prodt_end[57]) );
  CFD1QXL \prodt_end_reg[54]  ( .D(n262), .CP(clock), .Q(prodt_end[54]) );
  CFD1QXL \prodt_end_reg[53]  ( .D(n263), .CP(clock), .Q(prodt_end[53]) );
  CFD1QXL \prodt_end_reg[52]  ( .D(n264), .CP(clock), .Q(prodt_end[52]) );
  CFD1QXL \prodt_end_reg[60]  ( .D(n256), .CP(clock), .Q(prodt_end[60]) );
  CFD1QX1 \prodt_end_reg[48]  ( .D(n268), .CP(clock), .Q(prodt_end[48]) );
  CFD1QX1 \prodt_end_reg[49]  ( .D(n267), .CP(clock), .Q(prodt_end[49]) );
  CFD1QX1 \prodt_end_reg[55]  ( .D(n261), .CP(clock), .Q(prodt_end[55]) );
  CFD1QX1 \prodt_end_reg[47]  ( .D(n269), .CP(clock), .Q(prodt_end[47]) );
  CFD1QX1 \prodt_end_reg[50]  ( .D(n266), .CP(clock), .Q(prodt_end[50]) );
  CFD1QX1 \prodt_end_reg[56]  ( .D(n260), .CP(clock), .Q(prodt_end[56]) );
  CFD1QXL \prodt_end_reg[51]  ( .D(n265), .CP(clock), .Q(prodt_end[51]) );
  CFD1QXL \a_reg[31]  ( .D(n316), .CP(clock), .Q(a[31]) );
  CFD1QXL \a_reg[30]  ( .D(n317), .CP(clock), .Q(a[30]) );
  CFD1QXL \a_reg[29]  ( .D(n318), .CP(clock), .Q(a[29]) );
  CFD1QXL \a_reg[27]  ( .D(n320), .CP(clock), .Q(a[27]) );
  CFD1QXL \a_reg[23]  ( .D(n324), .CP(clock), .Q(a[23]) );
  CFD1QXL \a_reg[15]  ( .D(n332), .CP(clock), .Q(a[15]) );
  CFD1QXL \a_reg[28]  ( .D(n319), .CP(clock), .Q(a[28]) );
  CFD1QXL \a_reg[17]  ( .D(n330), .CP(clock), .Q(a[17]) );
  CFD1QXL \a_reg[12]  ( .D(n335), .CP(clock), .Q(a[12]) );
  CFD1QXL \a_reg[9]  ( .D(n338), .CP(clock), .Q(a[9]) );
  CFD1QXL \a_reg[10]  ( .D(n337), .CP(clock), .Q(a[10]) );
  CFD1QX1 \a_reg[5]  ( .D(n342), .CP(clock), .Q(a[5]) );
  CFD1QX1 \a_reg[8]  ( .D(n339), .CP(clock), .Q(a[8]) );
  CFD1QXL \prodt_end_reg[46]  ( .D(n270), .CP(clock), .Q(prodt_end[46]) );
  CFD1QXL \prodt_end_reg[43]  ( .D(n273), .CP(clock), .Q(prodt_end[43]) );
  CFD1QXL \prodt_end_reg[39]  ( .D(n277), .CP(clock), .Q(prodt_end[39]) );
  CFD1QXL \prodt_end_reg[45]  ( .D(n271), .CP(clock), .Q(prodt_end[45]) );
  CFD1QXL \prodt_end_reg[44]  ( .D(n272), .CP(clock), .Q(prodt_end[44]) );
  CFD1QXL \prodt_end_reg[42]  ( .D(n274), .CP(clock), .Q(prodt_end[42]) );
  CFD1QXL \prodt_end_reg[41]  ( .D(n275), .CP(clock), .Q(prodt_end[41]) );
  CFD1QXL \prodt_end_reg[38]  ( .D(n278), .CP(clock), .Q(prodt_end[38]) );
  CFD1QXL \prodt_end_reg[37]  ( .D(n279), .CP(clock), .Q(prodt_end[37]) );
  CFD1QXL \prodt_end_reg[35]  ( .D(n281), .CP(clock), .Q(prodt_end[35]) );
  CFD1QXL \prodt_end_reg[59]  ( .D(n257), .CP(clock), .Q(prodt_end[59]) );
  CFD1X1 \prodt_end_reg[40]  ( .D(n276), .CP(clock), .Q(prodt_end[40]), .QN(
        n419) );
  CFD1QX1 \a_reg[16]  ( .D(n331), .CP(clock), .Q(a[16]) );
  CFD1QX1 \a_reg[4]  ( .D(n343), .CP(clock), .Q(a[4]) );
  CFD1QX1 \a_reg[2]  ( .D(n345), .CP(clock), .Q(a[2]) );
  CFD1QX1 \prodt_end_reg[34]  ( .D(n282), .CP(clock), .Q(prodt_end[34]) );
  CFD1QX1 \prodt_end_reg[33]  ( .D(n283), .CP(clock), .Q(prodt_end[33]) );
  CFD1QX1 \prodt_end_reg[36]  ( .D(n280), .CP(clock), .Q(prodt_end[36]) );
  CFD1XL \count_reg[0]  ( .D(n412), .CP(clock), .Q(count[0]), .QN(n519) );
  CFD1QXL \a_reg[26]  ( .D(n321), .CP(clock), .Q(a[26]) );
  CFD1QXL \a_reg[25]  ( .D(n322), .CP(clock), .Q(a[25]) );
  CFD1QXL \a_reg[22]  ( .D(n325), .CP(clock), .Q(a[22]) );
  CFD1QXL \a_reg[21]  ( .D(n326), .CP(clock), .Q(a[21]) );
  CFD1QXL \a_reg[19]  ( .D(n328), .CP(clock), .Q(a[19]) );
  CFD1QXL \a_reg[14]  ( .D(n333), .CP(clock), .Q(a[14]) );
  CFD1QX1 \a_reg[13]  ( .D(n334), .CP(clock), .Q(a[13]) );
  CFD1QXL \a_reg[11]  ( .D(n336), .CP(clock), .Q(a[11]) );
  CFD1QXL \a_reg[7]  ( .D(n340), .CP(clock), .Q(a[7]) );
  CFD1QXL \a_reg[20]  ( .D(n327), .CP(clock), .Q(a[20]) );
  CFD1QXL \a_reg[18]  ( .D(n329), .CP(clock), .Q(a[18]) );
  CFD1QX1 \a_reg[1]  ( .D(n346), .CP(clock), .Q(a[1]) );
  CFD1QXL \a_reg[3]  ( .D(n344), .CP(clock), .Q(a[3]) );
  CFD1QXL \a_reg[6]  ( .D(n341), .CP(clock), .Q(a[6]) );
  CND2IX1 U405 ( .B(states[0]), .A(states[1]), .Z(n170) );
  CND2X1 U406 ( .A(count[5]), .B(n415), .Z(n522) );
  CENX1 U407 ( .A(mcand[0]), .B(a[0]), .Z(n215) );
  CND2X1 U408 ( .A(wsum[31]), .B(n424), .Z(n417) );
  CNR2X1 U409 ( .A(n459), .B(n164), .Z(n415) );
  CND2X1 U410 ( .A(prodt_end[63]), .B(n423), .Z(n416) );
  CAN2X1 U411 ( .A(n416), .B(n417), .Z(n97) );
  COND1X1 U412 ( .A(n427), .B(n450), .C(n104), .Z(n261) );
  COND1X1 U413 ( .A(n427), .B(n451), .C(n103), .Z(n260) );
  COND1X1 U414 ( .A(n427), .B(n442), .C(n112), .Z(n269) );
  COND1X1 U415 ( .A(n427), .B(n443), .C(n111), .Z(n268) );
  COND1X1 U416 ( .A(n427), .B(n444), .C(n110), .Z(n267) );
  COND1X1 U417 ( .A(n427), .B(n445), .C(n109), .Z(n266) );
  CIVX2 U418 ( .A(prodt_end[41]), .Z(n436) );
  CIVX2 U419 ( .A(prodt_end[42]), .Z(n437) );
  CIVX2 U420 ( .A(prodt_end[35]), .Z(n431) );
  CIVX2 U421 ( .A(prodt_end[38]), .Z(n434) );
  CIVX2 U422 ( .A(prodt_end[44]), .Z(n439) );
  CIVX1 U423 ( .A(prodt_end[51]), .Z(n446) );
  CANR2XL U424 ( .A(prodt_end[44]), .B(n422), .C(wsum[12]), .D(n96), .Z(n116)
         );
  CANR2XL U425 ( .A(prodt_end[45]), .B(n423), .C(wsum[13]), .D(n424), .Z(n115)
         );
  CANR2XL U426 ( .A(prodt_end[46]), .B(n95), .C(wsum[14]), .D(n424), .Z(n114)
         );
  CANR2XL U427 ( .A(prodt_end[40]), .B(n95), .C(wsum[8]), .D(n424), .Z(n120)
         );
  CANR2XL U428 ( .A(prodt_end[41]), .B(n422), .C(wsum[9]), .D(n424), .Z(n119)
         );
  CANR2XL U429 ( .A(prodt_end[42]), .B(n423), .C(wsum[10]), .D(n425), .Z(n118)
         );
  CANR2XL U430 ( .A(prodt_end[43]), .B(n95), .C(wsum[11]), .D(n425), .Z(n117)
         );
  CANR2XL U431 ( .A(prodt_end[36]), .B(n423), .C(wsum[4]), .D(n425), .Z(n124)
         );
  CANR2XL U432 ( .A(prodt_end[38]), .B(n422), .C(wsum[6]), .D(n96), .Z(n122)
         );
  CANR2XL U433 ( .A(prodt_end[39]), .B(n423), .C(wsum[7]), .D(n96), .Z(n121)
         );
  CANR2XL U434 ( .A(prodt_end[35]), .B(n422), .C(wsum[3]), .D(n425), .Z(n125)
         );
  CIVX2 U435 ( .A(prodt_end[37]), .Z(n433) );
  CAOR2XL U436 ( .A(n525), .B(a[1]), .C(n531), .D(mcand[1]), .Z(n346) );
  CAOR2XL U437 ( .A(n525), .B(a[10]), .C(n531), .D(mcand[10]), .Z(n337) );
  CAOR2XL U438 ( .A(n525), .B(a[5]), .C(n531), .D(mcand[5]), .Z(n342) );
  CAOR2XL U439 ( .A(n525), .B(a[8]), .C(n531), .D(mcand[8]), .Z(n339) );
  CAOR2XL U440 ( .A(n525), .B(a[3]), .C(n531), .D(mcand[3]), .Z(n344) );
  CAOR2XL U441 ( .A(n525), .B(a[6]), .C(n531), .D(mcand[6]), .Z(n341) );
  CIVX2 U442 ( .A(n131), .Z(n426) );
  CIVX2 U443 ( .A(n128), .Z(n532) );
  CIVX2 U444 ( .A(n415), .Z(n427) );
  CIVX2 U445 ( .A(n163), .Z(n531) );
  COND1XL U446 ( .A(n427), .B(n452), .C(n102), .Z(n259) );
  COND1XL U447 ( .A(n427), .B(n453), .C(n101), .Z(n258) );
  COND1XL U448 ( .A(n427), .B(n454), .C(n100), .Z(n257) );
  COND1XL U449 ( .A(n427), .B(n455), .C(n99), .Z(n256) );
  COND1XL U450 ( .A(n427), .B(n456), .C(n98), .Z(n255) );
  COND1XL U451 ( .A(n427), .B(n457), .C(n97), .Z(n254) );
  COND1XL U452 ( .A(n427), .B(n458), .C(n94), .Z(n253) );
  CND2X1 U453 ( .A(wcout), .B(n424), .Z(n94) );
  CND3XL U454 ( .A(n527), .B(n173), .C(n427), .Z(n128) );
  CAN8X1 U455 ( .A(n175), .B(n176), .C(n177), .D(n178), .E(n179), .F(n180), 
        .G(n181), .H(n182), .Z(n167) );
  CAN8X1 U456 ( .A(n241), .B(n242), .C(n243), .D(n244), .E(n245), .F(n246), 
        .G(n247), .H(n248), .Z(n175) );
  CAN8X1 U457 ( .A(n233), .B(n234), .C(n235), .D(n236), .E(n237), .F(n238), 
        .G(n239), .H(n240), .Z(n176) );
  CAN8X1 U458 ( .A(n225), .B(n226), .C(n227), .D(n228), .E(n229), .F(n230), 
        .G(n231), .H(n232), .Z(n177) );
  CND2X1 U459 ( .A(n527), .B(n526), .Z(n131) );
  CNR2X1 U460 ( .A(n537), .B(n131), .Z(n425) );
  CNR2X1 U461 ( .A(n537), .B(n131), .Z(n96) );
  CNR2X1 U462 ( .A(n537), .B(n131), .Z(n424) );
  CND2X1 U463 ( .A(n164), .B(n527), .Z(n163) );
  COND1XL U464 ( .A(n427), .B(n446), .C(n108), .Z(n265) );
  COND1XL U465 ( .A(n427), .B(n447), .C(n107), .Z(n264) );
  COND1XL U466 ( .A(n427), .B(n448), .C(n106), .Z(n263) );
  COND1XL U467 ( .A(n427), .B(n449), .C(n105), .Z(n262) );
  COND1XL U468 ( .A(n427), .B(n431), .C(n124), .Z(n281) );
  COND1XL U469 ( .A(n427), .B(n432), .C(n123), .Z(n280) );
  COND1XL U470 ( .A(n427), .B(n433), .C(n122), .Z(n279) );
  COND1XL U471 ( .A(n427), .B(n434), .C(n121), .Z(n278) );
  COND1XL U472 ( .A(n427), .B(n435), .C(n120), .Z(n277) );
  COND1XL U473 ( .A(n427), .B(n419), .C(n119), .Z(n276) );
  COND1XL U474 ( .A(n427), .B(n436), .C(n118), .Z(n275) );
  COND1XL U475 ( .A(n427), .B(n437), .C(n117), .Z(n274) );
  COND1XL U476 ( .A(n427), .B(n438), .C(n116), .Z(n273) );
  COND1XL U477 ( .A(n427), .B(n439), .C(n115), .Z(n272) );
  COND1XL U478 ( .A(n427), .B(n440), .C(n114), .Z(n271) );
  COND1XL U479 ( .A(n427), .B(n441), .C(n113), .Z(n270) );
  CANR2X1 U480 ( .A(prodt_end[47]), .B(n422), .C(wsum[15]), .D(n424), .Z(n113)
         );
  CIVX2 U481 ( .A(prodt_end[36]), .Z(n432) );
  CND2X1 U482 ( .A(prodt_end[31]), .B(n415), .Z(n129) );
  COND1XL U483 ( .A(n427), .B(n429), .C(n126), .Z(n283) );
  CANR2XL U484 ( .A(prodt_end[34]), .B(n95), .C(wsum[2]), .D(n425), .Z(n126)
         );
  COND1XL U485 ( .A(n427), .B(n430), .C(n125), .Z(n282) );
  CNR2X1 U486 ( .A(states[0]), .B(states[1]), .Z(n173) );
  CNR2X1 U487 ( .A(n534), .B(valid), .Z(n164) );
  COND1XL U488 ( .A(n427), .B(n567), .C(n172), .Z(n413) );
  CANR2X1 U489 ( .A(mlier[1]), .B(n532), .C(prodt_end[2]), .D(n426), .Z(n172)
         );
  COND1XL U490 ( .A(n427), .B(n566), .C(n160), .Z(n314) );
  CANR2X1 U491 ( .A(mlier[2]), .B(n532), .C(prodt_end[3]), .D(n426), .Z(n160)
         );
  COND1XL U492 ( .A(n427), .B(n565), .C(n159), .Z(n313) );
  CANR2X1 U493 ( .A(mlier[3]), .B(n532), .C(prodt_end[4]), .D(n426), .Z(n159)
         );
  COND1XL U494 ( .A(n427), .B(n564), .C(n158), .Z(n312) );
  CANR2X1 U495 ( .A(mlier[4]), .B(n532), .C(prodt_end[5]), .D(n426), .Z(n158)
         );
  COND1XL U496 ( .A(n427), .B(n563), .C(n157), .Z(n311) );
  CANR2X1 U497 ( .A(mlier[5]), .B(n532), .C(prodt_end[6]), .D(n426), .Z(n157)
         );
  COND1XL U498 ( .A(n427), .B(n562), .C(n156), .Z(n310) );
  CANR2X1 U499 ( .A(mlier[6]), .B(n532), .C(prodt_end[7]), .D(n426), .Z(n156)
         );
  COND1XL U500 ( .A(n427), .B(n561), .C(n155), .Z(n309) );
  CANR2X1 U501 ( .A(mlier[7]), .B(n532), .C(prodt_end[8]), .D(n426), .Z(n155)
         );
  COND1XL U502 ( .A(n427), .B(n560), .C(n154), .Z(n308) );
  CANR2X1 U503 ( .A(mlier[8]), .B(n532), .C(prodt_end[9]), .D(n426), .Z(n154)
         );
  COND1XL U504 ( .A(n427), .B(n559), .C(n153), .Z(n307) );
  CANR2X1 U505 ( .A(mlier[9]), .B(n532), .C(prodt_end[10]), .D(n426), .Z(n153)
         );
  COND1XL U506 ( .A(n427), .B(n558), .C(n152), .Z(n306) );
  CANR2X1 U507 ( .A(mlier[10]), .B(n532), .C(prodt_end[11]), .D(n426), .Z(n152) );
  COND1XL U508 ( .A(n427), .B(n557), .C(n151), .Z(n305) );
  CANR2X1 U509 ( .A(mlier[11]), .B(n532), .C(prodt_end[12]), .D(n426), .Z(n151) );
  COND1XL U510 ( .A(n427), .B(n556), .C(n150), .Z(n304) );
  CANR2X1 U511 ( .A(mlier[12]), .B(n532), .C(prodt_end[13]), .D(n426), .Z(n150) );
  COND1XL U512 ( .A(n427), .B(n555), .C(n149), .Z(n303) );
  CANR2X1 U513 ( .A(mlier[13]), .B(n532), .C(prodt_end[14]), .D(n426), .Z(n149) );
  COND1XL U514 ( .A(n427), .B(n554), .C(n148), .Z(n302) );
  CANR2X1 U515 ( .A(mlier[14]), .B(n532), .C(prodt_end[15]), .D(n426), .Z(n148) );
  COND1XL U516 ( .A(n427), .B(n553), .C(n147), .Z(n301) );
  CANR2X1 U517 ( .A(mlier[15]), .B(n532), .C(prodt_end[16]), .D(n426), .Z(n147) );
  COND1XL U518 ( .A(n427), .B(n552), .C(n146), .Z(n300) );
  CANR2X1 U519 ( .A(mlier[16]), .B(n532), .C(prodt_end[17]), .D(n426), .Z(n146) );
  COND1XL U520 ( .A(n427), .B(n551), .C(n145), .Z(n299) );
  CANR2X1 U521 ( .A(mlier[17]), .B(n532), .C(prodt_end[18]), .D(n426), .Z(n145) );
  COND1XL U522 ( .A(n427), .B(n550), .C(n144), .Z(n298) );
  CANR2X1 U523 ( .A(mlier[18]), .B(n532), .C(prodt_end[19]), .D(n426), .Z(n144) );
  COND1XL U524 ( .A(n427), .B(n549), .C(n143), .Z(n297) );
  CANR2X1 U525 ( .A(mlier[19]), .B(n532), .C(prodt_end[20]), .D(n426), .Z(n143) );
  COND1XL U526 ( .A(n427), .B(n548), .C(n142), .Z(n296) );
  CANR2X1 U527 ( .A(mlier[20]), .B(n532), .C(prodt_end[21]), .D(n426), .Z(n142) );
  COND1XL U528 ( .A(n427), .B(n547), .C(n141), .Z(n295) );
  CANR2X1 U529 ( .A(mlier[21]), .B(n532), .C(prodt_end[22]), .D(n426), .Z(n141) );
  COND1XL U530 ( .A(n427), .B(n546), .C(n140), .Z(n294) );
  CANR2X1 U531 ( .A(mlier[22]), .B(n532), .C(prodt_end[23]), .D(n426), .Z(n140) );
  COND1XL U532 ( .A(n427), .B(n545), .C(n139), .Z(n293) );
  CANR2X1 U533 ( .A(mlier[23]), .B(n532), .C(prodt_end[24]), .D(n426), .Z(n139) );
  COND1XL U534 ( .A(n427), .B(n544), .C(n138), .Z(n292) );
  CANR2X1 U535 ( .A(mlier[24]), .B(n532), .C(prodt_end[25]), .D(n426), .Z(n138) );
  COND1XL U536 ( .A(n427), .B(n543), .C(n137), .Z(n291) );
  CANR2X1 U537 ( .A(mlier[25]), .B(n532), .C(prodt_end[26]), .D(n426), .Z(n137) );
  COND1XL U538 ( .A(n427), .B(n542), .C(n136), .Z(n290) );
  CANR2X1 U539 ( .A(mlier[26]), .B(n532), .C(prodt_end[27]), .D(n426), .Z(n136) );
  COND1XL U540 ( .A(n427), .B(n541), .C(n135), .Z(n289) );
  CANR2X1 U541 ( .A(mlier[27]), .B(n532), .C(prodt_end[28]), .D(n426), .Z(n135) );
  COND1XL U542 ( .A(n427), .B(n540), .C(n134), .Z(n288) );
  CANR2X1 U543 ( .A(mlier[28]), .B(n532), .C(prodt_end[29]), .D(n426), .Z(n134) );
  COND1XL U544 ( .A(n427), .B(n539), .C(n133), .Z(n287) );
  CANR2X1 U545 ( .A(mlier[29]), .B(n532), .C(prodt_end[30]), .D(n426), .Z(n133) );
  COND1XL U546 ( .A(n427), .B(n538), .C(n132), .Z(n286) );
  CANR2X1 U547 ( .A(mlier[30]), .B(n532), .C(prodt_end[31]), .D(n426), .Z(n132) );
  CNR2IX1 U548 ( .B(count[30]), .A(n427), .Z(n461) );
  CNR2IX1 U549 ( .B(count[29]), .A(n427), .Z(n463) );
  CNR2IX1 U550 ( .B(count[28]), .A(n427), .Z(n465) );
  CNR2IX1 U551 ( .B(count[31]), .A(n427), .Z(n521) );
  COND2X1 U552 ( .A(n131), .B(n567), .C(n128), .D(n530), .Z(n161) );
  COND2X1 U553 ( .A(reset), .B(n534), .C(n535), .D(n131), .Z(N326) );
  CNR2X1 U554 ( .A(n131), .B(add), .Z(n422) );
  CNR2X1 U555 ( .A(n131), .B(add), .Z(n423) );
  CNR2X1 U556 ( .A(n131), .B(add), .Z(n95) );
  CENX1 U557 ( .A(mcand[4]), .B(a[4]), .Z(n210) );
  CENX1 U558 ( .A(mcand[3]), .B(a[3]), .Z(n209) );
  CENX1 U559 ( .A(mcand[2]), .B(a[2]), .Z(n208) );
  CENX1 U560 ( .A(mcand[1]), .B(a[1]), .Z(n207) );
  CND4X1 U561 ( .A(n249), .B(n250), .C(n251), .D(n252), .Z(n169) );
  COND2X1 U562 ( .A(n524), .B(n12), .C(n529), .D(n163), .Z(n348) );
  COND2X1 U563 ( .A(N326), .B(n537), .C(n533), .D(n174), .Z(n414) );
  CANR2X1 U564 ( .A(prodt_end[1]), .B(n526), .C(mlier[0]), .D(n173), .Z(n174)
         );
  CNR2X1 U565 ( .A(n223), .B(n224), .Z(n222) );
  CEOX1 U566 ( .A(mlier[27]), .B(b[27]), .Z(n223) );
  CEOX1 U567 ( .A(mlier[26]), .B(b[26]), .Z(n224) );
  CENX1 U568 ( .A(mcand[20]), .B(a[20]), .Z(n194) );
  CENX1 U569 ( .A(mcand[12]), .B(a[12]), .Z(n202) );
  CENX1 U570 ( .A(mcand[28]), .B(a[28]), .Z(n186) );
  CENX1 U571 ( .A(mlier[19]), .B(b[19]), .Z(n228) );
  CENX1 U572 ( .A(mlier[11]), .B(b[11]), .Z(n236) );
  CENX1 U573 ( .A(mlier[3]), .B(b[3]), .Z(n244) );
  CENX1 U574 ( .A(mcand[24]), .B(a[24]), .Z(n198) );
  CENX1 U575 ( .A(mcand[16]), .B(a[16]), .Z(n206) );
  CENX1 U576 ( .A(mcand[31]), .B(a[31]), .Z(n190) );
  CENX1 U577 ( .A(mlier[23]), .B(b[23]), .Z(n232) );
  CENX1 U578 ( .A(mlier[15]), .B(b[15]), .Z(n240) );
  CENX1 U579 ( .A(mlier[7]), .B(b[7]), .Z(n248) );
  CENX1 U580 ( .A(mcand[27]), .B(a[27]), .Z(n185) );
  CENX1 U581 ( .A(mlier[18]), .B(b[18]), .Z(n227) );
  CENX1 U582 ( .A(mlier[10]), .B(b[10]), .Z(n235) );
  CENX1 U583 ( .A(mlier[2]), .B(b[2]), .Z(n243) );
  CENX1 U584 ( .A(mlier[25]), .B(b[25]), .Z(n221) );
  CENX1 U585 ( .A(mcand[23]), .B(a[23]), .Z(n197) );
  CENX1 U586 ( .A(mcand[15]), .B(a[15]), .Z(n205) );
  CENX1 U587 ( .A(mlier[22]), .B(b[22]), .Z(n231) );
  CENX1 U588 ( .A(mlier[14]), .B(b[14]), .Z(n239) );
  CENX1 U589 ( .A(mlier[6]), .B(b[6]), .Z(n247) );
  CENX1 U590 ( .A(mlier[24]), .B(b[24]), .Z(n220) );
  CENX1 U591 ( .A(mcand[22]), .B(a[22]), .Z(n196) );
  CENX1 U592 ( .A(mcand[14]), .B(a[14]), .Z(n204) );
  CENX1 U593 ( .A(mcand[30]), .B(a[30]), .Z(n188) );
  CENX1 U594 ( .A(mlier[21]), .B(b[21]), .Z(n230) );
  CENX1 U595 ( .A(mlier[13]), .B(b[13]), .Z(n238) );
  CENX1 U596 ( .A(mlier[5]), .B(b[5]), .Z(n246) );
  CENX1 U597 ( .A(mcand[18]), .B(a[18]), .Z(n192) );
  CENX1 U598 ( .A(mlier[17]), .B(b[17]), .Z(n226) );
  CENX1 U599 ( .A(mlier[9]), .B(b[9]), .Z(n234) );
  CENX1 U600 ( .A(mlier[1]), .B(b[1]), .Z(n242) );
  CENX1 U601 ( .A(mlier[16]), .B(b[16]), .Z(n225) );
  CENX1 U602 ( .A(mlier[8]), .B(b[8]), .Z(n233) );
  CENX1 U603 ( .A(mlier[20]), .B(b[20]), .Z(n229) );
  CENX1 U604 ( .A(mlier[12]), .B(b[12]), .Z(n237) );
  CENX1 U605 ( .A(mlier[4]), .B(b[4]), .Z(n245) );
  COND1XL U606 ( .A(n427), .B(n511), .C(n510), .Z(n408) );
  COND1XL U607 ( .A(n427), .B(n513), .C(n512), .Z(n409) );
  CEOX1 U608 ( .A(mlier[31]), .B(n12), .Z(n217) );
  CEOX1 U609 ( .A(mlier[0]), .B(n13), .Z(n241) );
  COND1XL U610 ( .A(n427), .B(n519), .C(n518), .Z(n412) );
  CND2X1 U611 ( .A(N55), .B(n426), .Z(n518) );
  COND1XL U612 ( .A(n427), .B(n515), .C(n514), .Z(n410) );
  COND1XL U613 ( .A(n427), .B(n517), .C(n516), .Z(n411) );
  CND2X1 U614 ( .A(N56), .B(n426), .Z(n516) );
  COND1XL U615 ( .A(n165), .B(n536), .C(n166), .Z(n380) );
  COND3X1 U616 ( .A(n167), .B(n526), .C(n165), .D(n527), .Z(n166) );
  COND3X1 U617 ( .A(n528), .B(n169), .C(n527), .D(n170), .Z(n165) );
  CAN8X1 U618 ( .A(n215), .B(n216), .C(n217), .D(n218), .E(n219), .F(n220), 
        .G(n221), .H(n222), .Z(n178) );
  CENX1 U619 ( .A(mlier[29]), .B(b[29]), .Z(n219) );
  CENX1 U620 ( .A(mlier[30]), .B(b[30]), .Z(n216) );
  CENX1 U621 ( .A(mlier[28]), .B(b[28]), .Z(n218) );
  CAN8X1 U622 ( .A(n183), .B(n184), .C(n185), .D(n186), .E(n187), .F(n188), 
        .G(n189), .H(n190), .Z(n182) );
  CENX1 U623 ( .A(mcand[25]), .B(a[25]), .Z(n183) );
  CENX1 U624 ( .A(mcand[29]), .B(a[29]), .Z(n187) );
  CENX1 U625 ( .A(mcand[26]), .B(a[26]), .Z(n184) );
  CAN8X1 U626 ( .A(n191), .B(n192), .C(n193), .D(n194), .E(n195), .F(n196), 
        .G(n197), .H(n198), .Z(n181) );
  CENX1 U627 ( .A(mcand[17]), .B(a[17]), .Z(n191) );
  CENX1 U628 ( .A(mcand[21]), .B(a[21]), .Z(n195) );
  CENX1 U629 ( .A(mcand[19]), .B(a[19]), .Z(n193) );
  CAN8X1 U630 ( .A(n199), .B(n200), .C(n201), .D(n202), .E(n203), .F(n204), 
        .G(n205), .H(n206), .Z(n180) );
  CENX1 U631 ( .A(mcand[9]), .B(a[9]), .Z(n199) );
  CENX1 U632 ( .A(mcand[13]), .B(a[13]), .Z(n203) );
  CENX1 U633 ( .A(mcand[11]), .B(a[11]), .Z(n201) );
  CAN8X1 U634 ( .A(n207), .B(n208), .C(n209), .D(n210), .E(n211), .F(n212), 
        .G(n213), .H(n214), .Z(n179) );
  CENX1 U635 ( .A(mcand[7]), .B(a[7]), .Z(n213) );
  CENX1 U636 ( .A(mcand[8]), .B(a[8]), .Z(n214) );
  CND3XL U637 ( .A(n128), .B(n523), .C(n522), .Z(n407) );
  CNR2IX1 U638 ( .B(states[1]), .A(states[0]), .Z(n189) );
  CNR2IX1 U639 ( .B(count[27]), .A(n427), .Z(n467) );
  CNR2IX1 U640 ( .B(count[26]), .A(n427), .Z(n469) );
  CNR2IX1 U641 ( .B(count[25]), .A(n427), .Z(n471) );
  CNR2IX1 U642 ( .B(count[24]), .A(n427), .Z(n473) );
  CNR2IX1 U643 ( .B(count[23]), .A(n427), .Z(n475) );
  CNR2IX1 U644 ( .B(count[22]), .A(n427), .Z(n477) );
  CNR2IX1 U645 ( .B(count[21]), .A(n427), .Z(n479) );
  CNR2IX1 U646 ( .B(count[20]), .A(n427), .Z(n481) );
  CNR2IX1 U647 ( .B(count[19]), .A(n427), .Z(n483) );
  CNR2IX1 U648 ( .B(count[18]), .A(n427), .Z(n485) );
  CNR2IX1 U649 ( .B(count[17]), .A(n427), .Z(n487) );
  CNR2IX1 U650 ( .B(count[16]), .A(n427), .Z(n489) );
  CNR2IX1 U651 ( .B(count[15]), .A(n427), .Z(n491) );
  CNR2IX1 U652 ( .B(count[14]), .A(n427), .Z(n493) );
  CNR2IX1 U653 ( .B(count[13]), .A(n427), .Z(n495) );
  CNR2IX1 U654 ( .B(count[12]), .A(n427), .Z(n497) );
  CNR2IX1 U655 ( .B(count[11]), .A(n427), .Z(n499) );
  CNR2IX1 U656 ( .B(count[10]), .A(n427), .Z(n501) );
  CNR2IX1 U657 ( .B(count[9]), .A(n427), .Z(n503) );
  CNR2IX1 U658 ( .B(count[7]), .A(n427), .Z(n507) );
  COND2X1 U659 ( .A(n524), .B(n13), .C(n530), .D(n163), .Z(n379) );
  COND1XL U660 ( .A(n505), .B(n131), .C(n504), .Z(n404) );
  CND2X1 U661 ( .A(count[8]), .B(n415), .Z(n504) );
  COND1XL U662 ( .A(n509), .B(n131), .C(n508), .Z(n406) );
  CND2X1 U663 ( .A(count[6]), .B(n415), .Z(n508) );
  CAOR2XL U664 ( .A(n525), .B(a[0]), .C(n531), .D(mcand[0]), .Z(n347) );
  CIVXL U665 ( .A(prodt_end[32]), .Z(n428) );
  CANR2X1 U666 ( .A(prodt_end[48]), .B(n423), .C(wsum[16]), .D(n424), .Z(n112)
         );
  CANR2X1 U667 ( .A(prodt_end[55]), .B(n95), .C(wsum[23]), .D(n96), .Z(n105)
         );
  CANR2X1 U668 ( .A(prodt_end[54]), .B(n423), .C(wsum[22]), .D(n425), .Z(n106)
         );
  CANR2X1 U669 ( .A(prodt_end[53]), .B(n422), .C(wsum[21]), .D(n425), .Z(n107)
         );
  CANR2X1 U670 ( .A(prodt_end[52]), .B(n95), .C(wsum[20]), .D(n424), .Z(n108)
         );
  CANR2X1 U671 ( .A(prodt_end[51]), .B(n423), .C(wsum[19]), .D(n425), .Z(n109)
         );
  CANR2X1 U672 ( .A(prodt_end[50]), .B(n422), .C(wsum[18]), .D(n425), .Z(n110)
         );
  CANR2X1 U673 ( .A(prodt_end[49]), .B(n95), .C(wsum[17]), .D(n425), .Z(n111)
         );
  COND3X1 U674 ( .A(n128), .B(n529), .C(n129), .D(n130), .Z(n285) );
  CANR2XL U675 ( .A(prodt_end[32]), .B(n422), .C(wsum[0]), .D(n424), .Z(n130)
         );
  COND1XL U676 ( .A(n427), .B(n428), .C(n127), .Z(n284) );
  CIVX2 U677 ( .A(prodt_end[45]), .Z(n440) );
  CANR2X1 U678 ( .A(prodt_end[61]), .B(n95), .C(wsum[29]), .D(n424), .Z(n99)
         );
  CANR2X1 U679 ( .A(prodt_end[59]), .B(n422), .C(wsum[27]), .D(n96), .Z(n101)
         );
  CANR2X1 U680 ( .A(prodt_end[56]), .B(n422), .C(wsum[24]), .D(n425), .Z(n104)
         );
  CANR2X1 U681 ( .A(prodt_end[62]), .B(n422), .C(wsum[30]), .D(n424), .Z(n98)
         );
  CENX1 U682 ( .A(mcand[6]), .B(a[6]), .Z(n212) );
  CENX1 U683 ( .A(mcand[10]), .B(a[10]), .Z(n200) );
  CENX1 U684 ( .A(mcand[5]), .B(a[5]), .Z(n211) );
  CIVX2 U685 ( .A(prodt_end[56]), .Z(n451) );
  CANR2X1 U686 ( .A(prodt_end[60]), .B(n423), .C(wsum[28]), .D(n96), .Z(n100)
         );
  CIVX2 U687 ( .A(prodt_end[50]), .Z(n445) );
  CANR2X1 U688 ( .A(prodt_end[58]), .B(n95), .C(wsum[26]), .D(n96), .Z(n102)
         );
  CANR2X1 U689 ( .A(prodt_end[57]), .B(n423), .C(wsum[25]), .D(n96), .Z(n103)
         );
  CANR2XL U690 ( .A(prodt_end[37]), .B(n95), .C(wsum[5]), .D(n96), .Z(n123) );
  CAOR2XL U691 ( .A(n525), .B(a[2]), .C(n531), .D(mcand[2]), .Z(n345) );
  CANR2XL U692 ( .A(prodt_end[33]), .B(n423), .C(wsum[1]), .D(n425), .Z(n127)
         );
  CIVX1 U693 ( .A(prodt_end[33]), .Z(n429) );
  CIVX1 U694 ( .A(prodt_end[34]), .Z(n430) );
  CIVX1 U695 ( .A(prodt_end[39]), .Z(n435) );
  CIVX1 U696 ( .A(prodt_end[43]), .Z(n438) );
  CIVX1 U697 ( .A(prodt_end[46]), .Z(n441) );
  CIVX1 U698 ( .A(prodt_end[47]), .Z(n442) );
  CIVX1 U699 ( .A(prodt_end[48]), .Z(n443) );
  CIVX1 U700 ( .A(prodt_end[49]), .Z(n444) );
  CIVX1 U701 ( .A(prodt_end[52]), .Z(n447) );
  CIVX1 U702 ( .A(prodt_end[53]), .Z(n448) );
  CIVX1 U703 ( .A(prodt_end[54]), .Z(n449) );
  CIVX1 U704 ( .A(prodt_end[55]), .Z(n450) );
  CIVX1 U705 ( .A(prodt_end[57]), .Z(n452) );
  CIVX1 U706 ( .A(prodt_end[58]), .Z(n453) );
  CIVX1 U707 ( .A(prodt_end[59]), .Z(n454) );
  CIVX1 U708 ( .A(prodt_end[60]), .Z(n455) );
  CIVX1 U709 ( .A(prodt_end[61]), .Z(n456) );
  CIVX1 U710 ( .A(prodt_end[62]), .Z(n457) );
  CIVX1 U711 ( .A(prodt_end[63]), .Z(n458) );
  CND2IX1 U712 ( .B(states[1]), .A(states[0]), .Z(n528) );
  CND2IX1 U713 ( .B(reset), .A(n528), .Z(n459) );
  CIVX2 U714 ( .A(reset), .Z(n527) );
  CIVX2 U715 ( .A(n528), .Z(n526) );
  CND2IX1 U716 ( .B(n131), .A(N85), .Z(n460) );
  CND2IX1 U717 ( .B(n461), .A(n460), .Z(n382) );
  CND2IX1 U718 ( .B(n131), .A(N84), .Z(n462) );
  CND2IX1 U719 ( .B(n463), .A(n462), .Z(n383) );
  CND2IX1 U720 ( .B(n131), .A(N83), .Z(n464) );
  CND2IX1 U721 ( .B(n465), .A(n464), .Z(n384) );
  CND2IX1 U722 ( .B(n131), .A(N82), .Z(n466) );
  CND2IX1 U723 ( .B(n467), .A(n466), .Z(n385) );
  CND2IX1 U724 ( .B(n131), .A(N81), .Z(n468) );
  CND2IX1 U725 ( .B(n469), .A(n468), .Z(n386) );
  CND2IX1 U726 ( .B(n131), .A(N80), .Z(n470) );
  CND2IX1 U727 ( .B(n471), .A(n470), .Z(n387) );
  CND2IX1 U728 ( .B(n131), .A(N79), .Z(n472) );
  CND2IX1 U729 ( .B(n473), .A(n472), .Z(n388) );
  CND2IX1 U730 ( .B(n131), .A(N78), .Z(n474) );
  CND2IX1 U731 ( .B(n475), .A(n474), .Z(n389) );
  CND2IX1 U732 ( .B(n131), .A(N77), .Z(n476) );
  CND2IX1 U733 ( .B(n477), .A(n476), .Z(n390) );
  CND2IX1 U734 ( .B(n131), .A(N76), .Z(n478) );
  CND2IX1 U735 ( .B(n479), .A(n478), .Z(n391) );
  CND2IX1 U736 ( .B(n131), .A(N75), .Z(n480) );
  CND2IX1 U737 ( .B(n481), .A(n480), .Z(n392) );
  CND2IX1 U738 ( .B(n131), .A(N74), .Z(n482) );
  CND2IX1 U739 ( .B(n483), .A(n482), .Z(n393) );
  CND2IX1 U740 ( .B(n131), .A(N73), .Z(n484) );
  CND2IX1 U741 ( .B(n485), .A(n484), .Z(n394) );
  CND2IX1 U742 ( .B(n131), .A(N72), .Z(n486) );
  CND2IX1 U743 ( .B(n487), .A(n486), .Z(n395) );
  CND2IX1 U744 ( .B(n131), .A(N71), .Z(n488) );
  CND2IX1 U745 ( .B(n489), .A(n488), .Z(n396) );
  CND2IX1 U746 ( .B(n131), .A(N70), .Z(n490) );
  CND2IX1 U747 ( .B(n491), .A(n490), .Z(n397) );
  CND2IX1 U748 ( .B(n131), .A(N69), .Z(n492) );
  CND2IX1 U749 ( .B(n493), .A(n492), .Z(n398) );
  CND2IX1 U750 ( .B(n131), .A(N68), .Z(n494) );
  CND2IX1 U751 ( .B(n495), .A(n494), .Z(n399) );
  CND2IX1 U752 ( .B(n131), .A(N67), .Z(n496) );
  CND2IX1 U753 ( .B(n497), .A(n496), .Z(n400) );
  CND2IX1 U754 ( .B(n131), .A(N66), .Z(n498) );
  CND2IX1 U755 ( .B(n499), .A(n498), .Z(n401) );
  CND2IX1 U756 ( .B(n131), .A(N65), .Z(n500) );
  CND2IX1 U757 ( .B(n501), .A(n500), .Z(n402) );
  CND2IX1 U758 ( .B(n131), .A(N64), .Z(n502) );
  CND2IX1 U759 ( .B(n503), .A(n502), .Z(n403) );
  CIVX2 U760 ( .A(N63), .Z(n505) );
  CND2IX1 U761 ( .B(n131), .A(N62), .Z(n506) );
  CND2IX1 U762 ( .B(n507), .A(n506), .Z(n405) );
  CIVX2 U763 ( .A(N61), .Z(n509) );
  CIVX2 U764 ( .A(count[4]), .Z(n511) );
  CND2IX1 U765 ( .B(n131), .A(N59), .Z(n510) );
  CIVX2 U766 ( .A(count[3]), .Z(n513) );
  CND2IX1 U767 ( .B(n131), .A(N58), .Z(n512) );
  CIVX2 U768 ( .A(count[2]), .Z(n515) );
  CND2IX1 U769 ( .B(n131), .A(N57), .Z(n514) );
  CIVX2 U770 ( .A(count[1]), .Z(n517) );
  CND2IX1 U771 ( .B(n131), .A(N86), .Z(n520) );
  CND2IX1 U772 ( .B(n521), .A(n520), .Z(n381) );
  CND2IX1 U773 ( .B(n131), .A(N60), .Z(n523) );
  CND2IX1 U774 ( .B(n164), .A(n527), .Z(n524) );
  CIVX2 U775 ( .A(n524), .Z(n525) );
  CIVX2 U776 ( .A(mlier[31]), .Z(n529) );
  CIVX2 U777 ( .A(mlier[0]), .Z(n530) );
  CIVX2 U778 ( .A(N326), .Z(n533) );
  CIVX2 U779 ( .A(n173), .Z(n534) );
  CIVX2 U780 ( .A(n169), .Z(n535) );
  CIVX2 U781 ( .A(valid), .Z(n536) );
  CIVX2 U782 ( .A(add), .Z(n537) );
  CIVX2 U783 ( .A(prodt_end[30]), .Z(n538) );
  CIVX2 U784 ( .A(prodt_end[29]), .Z(n539) );
  CIVX2 U785 ( .A(prodt_end[28]), .Z(n540) );
  CIVX2 U786 ( .A(prodt_end[27]), .Z(n541) );
  CIVX2 U787 ( .A(prodt_end[26]), .Z(n542) );
  CIVX2 U788 ( .A(prodt_end[25]), .Z(n543) );
  CIVX2 U789 ( .A(prodt_end[24]), .Z(n544) );
  CIVX2 U790 ( .A(prodt_end[23]), .Z(n545) );
  CIVX2 U791 ( .A(prodt_end[22]), .Z(n546) );
  CIVX2 U792 ( .A(prodt_end[21]), .Z(n547) );
  CIVX2 U793 ( .A(prodt_end[20]), .Z(n548) );
  CIVX2 U794 ( .A(prodt_end[19]), .Z(n549) );
  CIVX2 U795 ( .A(prodt_end[18]), .Z(n550) );
  CIVX2 U796 ( .A(prodt_end[17]), .Z(n551) );
  CIVX2 U797 ( .A(prodt_end[16]), .Z(n552) );
  CIVX2 U798 ( .A(prodt_end[15]), .Z(n553) );
  CIVX2 U799 ( .A(prodt_end[14]), .Z(n554) );
  CIVX2 U800 ( .A(prodt_end[13]), .Z(n555) );
  CIVX2 U801 ( .A(prodt_end[12]), .Z(n556) );
  CIVX2 U802 ( .A(prodt_end[11]), .Z(n557) );
  CIVX2 U803 ( .A(prodt_end[10]), .Z(n558) );
  CIVX2 U804 ( .A(prodt_end[9]), .Z(n559) );
  CIVX2 U805 ( .A(prodt_end[8]), .Z(n560) );
  CIVX2 U806 ( .A(prodt_end[7]), .Z(n561) );
  CIVX2 U807 ( .A(prodt_end[6]), .Z(n562) );
  CIVX2 U808 ( .A(prodt_end[5]), .Z(n563) );
  CIVX2 U809 ( .A(prodt_end[4]), .Z(n564) );
  CIVX2 U810 ( .A(prodt_end[3]), .Z(n565) );
  CIVX2 U811 ( .A(prodt_end[2]), .Z(n566) );
  CIVX2 U812 ( .A(prodt_end[1]), .Z(n567) );
endmodule

