
module Add_half_0 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7679 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_0 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_0 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7679 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_7673 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7674 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX2 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3837 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7674 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7673 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7675 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7676 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX2 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3838 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7676 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7675 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7677 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7678 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3839 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7678 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7677 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_0 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_0 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0)
         );
  Add_full_3839 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3838 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3837 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s3), .Z(n5) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CANR2X4 U5 ( .A(n1), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n4) );
  CIVX2 U6 ( .A(c_out11), .Z(n3) );
  CIVX2 U7 ( .A(c_out10), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n6) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_7649 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7650 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3825 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7650 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7649 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7651 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7652 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3826 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7652 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7651 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7653 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7654 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3827 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7654 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7653 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_7655 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7656 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3828 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7656 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7655 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_957 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3828 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3827 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3826 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3825 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_7657 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7658 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3829 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7658 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7657 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7659 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7660 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3830 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7660 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7659 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7661 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7662 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3831 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7662 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7661 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_7663 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7664 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3832 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7664 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7663 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_958 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3832 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3831 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3830 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3829 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_7665 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7666 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX2 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3833 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7666 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7665 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_7667 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
  CIVX2 U4 ( .A(b), .Z(n2) );
endmodule


module Add_half_7668 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX2 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3834 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7668 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7667 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_7669 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7670 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net87622, n1;
  assign c_out = net87622;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(net87622) );
endmodule


module Add_full_3835 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7670 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7669 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n1), .B(n2), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n2) );
  CIVX2 U3 ( .A(w3), .Z(n1) );
endmodule


module Add_half_7671 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7672 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3836 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7672 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7671 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_959 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, net91982,
         net84743, net84742, n1, n2, n3, n4;

  Add_full_3836 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3835 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3834 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3833 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2X1 U3 ( .A(n4), .B(c_out00), .Z(n2) );
  CND2X2 U4 ( .A(c_in2), .B(c_out01), .Z(n3) );
  CND2X2 U5 ( .A(n2), .B(n3), .Z(n1) );
  CMXI2X1 U6 ( .A0(net84743), .A1(net84742), .S(n1), .Z(c_out2) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMX2X1 U8 ( .A0(s4), .A1(s3), .S(net91982), .Z(sum2[1]) );
  CIVX2 U9 ( .A(c_in2), .Z(n4) );
  CANR2X1 U10 ( .A(n4), .B(c_out00), .C(c_in2), .D(c_out01), .Z(net91982) );
  CIVX2 U11 ( .A(c_out10), .Z(net84743) );
  CIVX2 U12 ( .A(c_out11), .Z(net84742) );
endmodule


module bit4_0 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, net84778, net84779, net84782,
         net84783, net84785, net84784, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_0 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_959 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_958 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_957 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(n6), .A1(n5), .S(n1), .Z(sum4[3]) );
  CANR2XL U4 ( .A(n4), .B(c_out400), .C(c_in4), .D(c_out401), .Z(n1) );
  CANR2XL U5 ( .A(n4), .B(c_out400), .C(c_in4), .D(c_out401), .Z(n2) );
  CMXI2X1 U6 ( .A0(net84784), .A1(net84785), .S(n3), .Z(c_out4) );
  CIVX2 U7 ( .A(c_out410), .Z(net84785) );
  CIVX2 U8 ( .A(c_out411), .Z(net84784) );
  CANR2X1 U9 ( .A(n4), .B(c_out400), .C(c_in4), .D(c_out401), .Z(n3) );
  CMXI2XL U10 ( .A0(net84778), .A1(net84779), .S(n2), .Z(sum4[2]) );
  CIVX2 U11 ( .A(c_in4), .Z(n4) );
  CMXI2X1 U12 ( .A0(net84782), .A1(net84783), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U13 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX1 U14 ( .A(s42[0]), .Z(net84783) );
  CIVX1 U15 ( .A(s41[0]), .Z(net84782) );
  CIVX2 U16 ( .A(s44[0]), .Z(net84778) );
  CIVX2 U17 ( .A(s43[0]), .Z(net84779) );
  CIVX2 U18 ( .A(s44[1]), .Z(n6) );
  CIVX2 U19 ( .A(s43[1]), .Z(n5) );
endmodule


module Add_half_7553 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7554 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3777 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7554 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7553 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7555 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7556 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3778 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7556 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7555 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7557 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7558 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3779 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7558 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7557 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7559 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7560 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3780 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7560 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7559 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_945 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3780 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3779 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3778 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3777 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_7561 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7562 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3781 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7562 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7561 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7563 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7564 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3782 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7564 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7563 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7565 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7566 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3783 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7566 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7565 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7567 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7568 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3784 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7568 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7567 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_946 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_3784 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3783 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3782 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3781 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_7569 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7570 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3785 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7570 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7569 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7571 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7572 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3786 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7572 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7571 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7573 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7574 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3787 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7574 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7573 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7575 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7576 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3788 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7576 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7575 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_947 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3788 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3787 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3786 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3785 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n3) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVXL U6 ( .A(n2), .Z(n6) );
  CMXI2X1 U7 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CMX2XL U8 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CMX2X1 U9 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U10 ( .A(c_out10), .Z(n5) );
  CIVX2 U11 ( .A(c_out11), .Z(n4) );
endmodule


module Add_half_7577 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7578 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3789 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7578 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7577 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7579 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7580 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3790 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7580 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7579 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7581 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7582 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3791 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7582 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7581 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7583 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7584 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3792 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7584 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7583 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_948 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3792 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3791 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3790 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3789 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMX2XL U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U5 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out10), .Z(n4) );
  CIVX2 U9 ( .A(c_out11), .Z(n3) );
endmodule


module bit4_237 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_948 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_947 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_946 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_945 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n9), .A1(n8), .S(n1), .Z(sum4[3]) );
  CMXI2XL U4 ( .A0(n7), .A1(n6), .S(n1), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CMX2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(s41[0]), .Z(n3) );
  CIVX2 U8 ( .A(s42[0]), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U10 ( .A(s41[1]), .Z(n5) );
  CIVX2 U11 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U13 ( .A(s43[0]), .Z(n7) );
  CIVX2 U14 ( .A(s44[0]), .Z(n6) );
  CIVX2 U15 ( .A(s43[1]), .Z(n9) );
  CIVX2 U16 ( .A(s44[1]), .Z(n8) );
endmodule


module Add_half_7585 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7586 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3793 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7586 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7585 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7587 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7588 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3794 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7588 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7587 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7589 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7590 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3795 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7590 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7589 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7591 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7592 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVXL U1 ( .A(a), .Z(n1) );
  CENXL U2 ( .A(n1), .B(b), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3796 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7592 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7591 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_949 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_3796 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3795 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3794 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3793 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_7593 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7594 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3797 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7594 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7593 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7595 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7596 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3798 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7596 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7595 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7597 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7598 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3799 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7598 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7597 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7599 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7600 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3800 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7600 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7599 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_950 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_3800 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3799 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3798 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3797 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_7601 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7602 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3801 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7602 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7601 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7603 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7604 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3802 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7604 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7603 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7605 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7606 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3803 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7606 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7605 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7607 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7608 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3804 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7608 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7607 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_951 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n2, n3, n4, n5,
         n6, n7, n8, n9;

  Add_full_3804 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3803 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3802 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3801 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CIVDXL U4 ( .A(n2), .Z0(n7) );
  CIVX2 U5 ( .A(c_out10), .Z(n4) );
  CIVX2 U6 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX2 U8 ( .A(s1), .Z(n6) );
  CIVX2 U9 ( .A(s2), .Z(n5) );
  CMXI2X1 U10 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n9) );
  CIVX2 U12 ( .A(s4), .Z(n8) );
  CMXI2X1 U13 ( .A0(n9), .A1(n8), .S(n7), .Z(sum2[1]) );
endmodule


module Add_half_7609 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7610 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3805 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7610 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7609 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7611 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7612 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3806 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7612 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7611 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7613 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_7614 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3807 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7614 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7613 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7615 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7616 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3808 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7616 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7615 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_952 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3808 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3807 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3806 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3805 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMX2XL U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n4) );
  CIVX2 U8 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module bit4_238 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_952 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_951 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_950 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_949 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(c_in4), .Z(n1) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n2), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(c_out401), .A1(c_out400), .S(n1), .Z(n2) );
  CMX2XL U6 ( .A0(s43[1]), .A1(s44[1]), .S(n2), .Z(sum4[3]) );
  CMX2X1 U7 ( .A0(c_out410), .A1(c_out411), .S(n3), .Z(c_out4) );
  CMX2X1 U8 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U9 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n3) );
endmodule


module Add_half_7617 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_7618 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3809 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7618 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7617 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7619 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7620 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3810 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7620 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7619 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7621 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7622 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3811 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7622 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7621 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_7623 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7624 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3812 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7624 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7623 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_953 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_3812 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3811 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3810 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3809 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n7), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_out10), .Z(n4) );
  CIVX2 U7 ( .A(c_out11), .Z(n3) );
  CIVX2 U8 ( .A(n2), .Z(n7) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n7), .Z(c_out2) );
  CIVX2 U10 ( .A(s1), .Z(n6) );
  CIVX2 U11 ( .A(s2), .Z(n5) );
  CMXI2X1 U12 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_7625 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7626 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3813 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7626 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7625 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7627 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7628 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3814 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7628 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7627 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7629 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CENX1 U4 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7630 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3815 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7630 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7629 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7631 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(n1), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
  CND2X1 U3 ( .A(a), .B(b), .Z(n1) );
endmodule


module Add_half_7632 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3816 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7632 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7631 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_954 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3816 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3815 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3814 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3813 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s4), .Z(n5) );
  CIVX1 U4 ( .A(s3), .Z(n6) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n4) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_7633 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7634 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX2 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3817 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7634 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7633 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_7635 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3;

  CEOX1 U1 ( .A(n1), .B(n3), .Z(sum) );
  CIVX1 U2 ( .A(a), .Z(n1) );
  CND2X2 U3 ( .A(a), .B(b), .Z(n2) );
  CIVX2 U4 ( .A(n2), .Z(c_out) );
  CIVX2 U5 ( .A(b), .Z(n3) );
endmodule


module Add_half_7636 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX4 U1 ( .A(a), .Z(n1) );
  CENX2 U2 ( .A(n1), .B(b), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3818 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7636 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7635 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_7637 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CNIVX2 U1 ( .A(a), .Z(n2) );
  CND2X2 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
  CEOX2 U4 ( .A(b), .B(n2), .Z(sum) );
endmodule


module Add_half_7638 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net87621, n1;
  assign c_out = net87621;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX2 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(net87621) );
endmodule


module Add_full_3819 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7638 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7637 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n1), .B(n2), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n2) );
  CIVX2 U3 ( .A(w3), .Z(n1) );
endmodule


module Add_half_7639 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n3;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(n1), .B(a), .Z(sum) );
  CND2X2 U3 ( .A(a), .B(b), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(c_out) );
endmodule


module Add_half_7640 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(n1), .B(a), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3820 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7640 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7639 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_955 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, net84612,
         net84613, net91018, net84615, net84614, n1, n2, n3, n4;

  Add_full_3820 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3819 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3818 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3817 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(s2), .Z(net84613) );
  CND2X2 U4 ( .A(c_out00), .B(n4), .Z(n2) );
  CND2X1 U5 ( .A(c_in2), .B(c_out01), .Z(n3) );
  CND2X2 U6 ( .A(n2), .B(n3), .Z(n1) );
  CMXI2X1 U7 ( .A0(net84615), .A1(net84614), .S(n1), .Z(c_out2) );
  CIVX2 U8 ( .A(c_in2), .Z(n4) );
  CANR2X1 U9 ( .A(c_out00), .B(n4), .C(c_in2), .D(c_out01), .Z(net91018) );
  CIVX2 U10 ( .A(c_out10), .Z(net84615) );
  CIVX2 U11 ( .A(c_out11), .Z(net84614) );
  CMXI2X1 U12 ( .A0(net84612), .A1(net84613), .S(c_in2), .Z(sum2[0]) );
  CIVX1 U13 ( .A(s1), .Z(net84612) );
  CMX2X1 U14 ( .A0(s4), .A1(s3), .S(net91018), .Z(sum2[1]) );
endmodule


module Add_half_7641 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7642 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX2 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3821 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7642 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7641 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7643 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
  CIVX2 U4 ( .A(b), .Z(n2) );
endmodule


module Add_half_7644 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX2 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3822 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7644 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7643 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7645 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVX2 U1 ( .A(n1), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CND2X1 U3 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U4 ( .A(b), .Z(n2) );
endmodule


module Add_half_7646 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3823 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7646 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7645 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_7647 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
  CND2X1 U3 ( .A(a), .B(b), .Z(n1) );
endmodule


module Add_half_7648 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3824 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7648 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7647 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_956 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_3824 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3823 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3822 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3821 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s4), .A1(s3), .S(n5), .Z(sum2[1]) );
  CANR2X2 U4 ( .A(n2), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n1) );
  CANR2X1 U5 ( .A(n2), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n5) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out11), .Z(n4) );
  CIVX2 U8 ( .A(c_out10), .Z(n3) );
  CIVX2 U9 ( .A(c_in2), .Z(n2) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(n1), .Z(c_out2) );
endmodule


module bit4_239 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, net89861, net89860, net84657,
         net84656, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_956 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_955 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_954 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_953 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out400), .B(n2), .C(c_in4), .D(c_out401), .Z(n1) );
  CMXI2X1 U4 ( .A0(net84656), .A1(net84657), .S(n1), .Z(c_out4) );
  CIVXL U5 ( .A(n1), .Z(net89860) );
  CIVX2 U6 ( .A(c_in4), .Z(n2) );
  CMX2X1 U7 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U8 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX1 U9 ( .A(c_out410), .Z(net84657) );
  CIVX1 U10 ( .A(c_out411), .Z(net84656) );
  CIVX2 U11 ( .A(net89860), .Z(net89861) );
  CMXI2X1 U12 ( .A0(n4), .A1(n3), .S(net89861), .Z(sum4[2]) );
  CMXI2XL U13 ( .A0(n6), .A1(n5), .S(net89861), .Z(sum4[3]) );
  CIVX2 U14 ( .A(s44[0]), .Z(n4) );
  CIVX2 U15 ( .A(s43[0]), .Z(n3) );
  CIVX2 U16 ( .A(s44[1]), .Z(n6) );
  CIVX2 U17 ( .A(s43[1]), .Z(n5) );
endmodule


module bit8_0 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   n9, n10, c_out800, c_out801, c_out810, c_out811, net84790, net84791,
         net84800, net89758, net91652, net91898, net84795, net84794, net108263,
         net90142, net84806, net84805, net84789, n1, n3, n4, n5, n6, n7, n8;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;
  assign sum8[6] = net89758;

  bit4_0 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4({b8[3:2], n1, 
        b8[0]}), .c_in4(1'b0) );
  bit4_239 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4({b8[3:2], n4, 
        b8[0]}), .c_in4(1'b1) );
  bit4_238 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_237 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVX2 U3 ( .A(c_in8), .Z(net91898) );
  CIVX8 U4 ( .A(n3), .Z(n1) );
  CIVX8 U5 ( .A(n3), .Z(n4) );
  CMXI2X1 U6 ( .A0(net84805), .A1(net84806), .S(net84789), .Z(c_out8) );
  CANR2X1 U7 ( .A(c_out800), .B(net84800), .C(c_in8), .D(c_out801), .Z(
        net84789) );
  CANR2X1 U8 ( .A(c_out800), .B(net84800), .C(c_in8), .D(c_out801), .Z(
        net91652) );
  CANR2X1 U9 ( .A(c_out800), .B(net84800), .C(c_in8), .D(c_out801), .Z(
        net90142) );
  CIVX1 U10 ( .A(c_out810), .Z(net84806) );
  CIVX2 U11 ( .A(c_out811), .Z(net84805) );
  CMXI2X1 U12 ( .A0(net84794), .A1(net84795), .S(net90142), .Z(sum8[4]) );
  CMXI2XL U13 ( .A0(net84790), .A1(net84791), .S(net90142), .Z(n9) );
  CNIVX4 U14 ( .A(n10), .Z(sum8[0]) );
  CMX2X1 U15 ( .A0(s82[0]), .A1(s81[0]), .S(net91898), .Z(n10) );
  CMX2X1 U16 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CNIVX1 U17 ( .A(net91652), .Z(net108263) );
  CIVX2 U18 ( .A(s83[0]), .Z(net84795) );
  CIVX2 U19 ( .A(s84[0]), .Z(net84794) );
  CMX2X1 U20 ( .A0(s84[3]), .A1(s83[3]), .S(net108263), .Z(sum8[7]) );
  CIVXL U21 ( .A(s84[2]), .Z(net84790) );
  CIVX4 U22 ( .A(b8[1]), .Z(n3) );
  CMX2X2 U23 ( .A0(s84[1]), .A1(s83[1]), .S(net91652), .Z(sum8[5]) );
  CIVXL U24 ( .A(s83[2]), .Z(net84791) );
  CND2X4 U25 ( .A(n8), .B(n7), .Z(sum8[2]) );
  CND2IX2 U26 ( .B(net84800), .A(s82[2]), .Z(n7) );
  CNIVX3 U27 ( .A(n9), .Z(net89758) );
  CIVX2 U28 ( .A(s81[1]), .Z(n6) );
  CIVX2 U29 ( .A(s82[1]), .Z(n5) );
  CMXI2X1 U30 ( .A0(n6), .A1(n5), .S(c_in8), .Z(sum8[1]) );
  CND2IX1 U31 ( .B(c_in8), .A(s81[2]), .Z(n8) );
  CIVX2 U32 ( .A(c_in8), .Z(net84800) );
endmodule


module Add_half_7169 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7170 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3585 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7170 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7169 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7171 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7172 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3586 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7172 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7171 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7173 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7174 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3587 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7174 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7173 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7175 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7176 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3588 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7176 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7175 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_897 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3588 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3587 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3586 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3585 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7177 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7178 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3589 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7178 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7177 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7179 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7180 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3590 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7180 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7179 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7181 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7182 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3591 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7182 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7181 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7183 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7184 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3592 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7184 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7183 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_898 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3592 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3591 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3590 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3589 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7185 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7186 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3593 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7186 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7185 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7187 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7188 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3594 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7188 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7187 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7189 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7190 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3595 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7190 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7189 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7191 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7192 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3596 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7192 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7191 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_899 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3596 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3595 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3594 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3593 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7193 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7194 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3597 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7194 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7193 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7195 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7196 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3598 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7196 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7195 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7197 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7198 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3599 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7198 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7197 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7199 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7200 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3600 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7200 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7199 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_900 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3600 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3599 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3598 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3597 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_225 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_900 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_899 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_898 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_897 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_7201 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7202 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3601 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7202 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7201 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7203 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7204 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3602 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7204 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7203 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7205 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7206 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3603 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7206 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7205 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7207 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7208 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3604 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7208 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7207 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_901 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3604 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3603 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3602 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3601 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7209 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7210 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3605 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7210 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7209 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7211 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7212 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3606 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7212 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7211 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7213 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7214 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3607 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7214 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7213 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7215 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7216 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3608 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7216 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7215 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_902 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3608 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3607 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3606 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3605 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7217 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7218 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3609 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7218 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7217 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7219 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7220 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3610 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7220 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7219 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7221 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7222 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3611 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7222 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7221 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7223 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7224 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3612 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7224 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7223 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_903 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3612 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3611 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3610 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3609 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7225 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7226 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3613 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7226 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7225 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7227 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7228 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3614 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7228 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7227 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7229 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7230 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3615 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7230 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7229 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7231 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7232 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3616 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7232 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7231 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_904 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3616 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3615 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3614 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3613 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_226 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_904 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_903 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_902 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_901 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_7233 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7234 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3617 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7234 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7233 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7235 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7236 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3618 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7236 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7235 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7237 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7238 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3619 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7238 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7237 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7239 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7240 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3620 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7240 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7239 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_905 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3620 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3619 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3618 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3617 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7241 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7242 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3621 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7242 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7241 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7243 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7244 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3622 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7244 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7243 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7245 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7246 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3623 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7246 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7245 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7247 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7248 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3624 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7248 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7247 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_906 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3624 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3623 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3622 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3621 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7249 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7250 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3625 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7250 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7249 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7251 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7252 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3626 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7252 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7251 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7253 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7254 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3627 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7254 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7253 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7255 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7256 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3628 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7256 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7255 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_907 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3628 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3627 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3626 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3625 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7257 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7258 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3629 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7258 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7257 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7259 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7260 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3630 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7260 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7259 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7261 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7262 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3631 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7262 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7261 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7263 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7264 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3632 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7264 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7263 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_908 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3632 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3631 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3630 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3629 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_227 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_908 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_907 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_906 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_905 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_7265 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7266 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3633 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7266 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7265 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7267 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7268 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3634 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7268 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7267 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7269 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7270 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3635 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7270 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7269 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7271 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7272 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3636 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7272 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7271 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_909 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3636 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3635 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3634 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3633 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7273 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7274 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3637 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7274 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7273 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7275 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7276 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3638 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7276 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7275 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7277 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7278 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3639 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7278 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7277 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7279 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7280 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3640 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7280 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7279 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_910 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3640 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3639 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3638 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3637 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7281 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7282 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3641 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7282 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7281 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7283 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7284 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3642 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7284 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7283 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7285 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7286 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3643 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7286 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7285 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7287 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7288 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3644 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7288 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7287 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_911 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3644 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3643 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3642 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3641 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7289 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7290 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3645 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7290 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7289 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7291 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7292 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3646 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7292 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7291 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7293 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7294 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3647 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7294 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7293 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7295 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7296 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3648 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7296 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7295 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_912 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3648 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3647 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3646 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3645 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_228 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_912 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_911 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_910 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_909 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_57 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_228 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_227 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_226 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_225 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMXI2X2 U3 ( .A0(n2), .A1(n3), .S(n4), .Z(sum8[3]) );
  CIVX2 U4 ( .A(s81[3]), .Z(n2) );
  CIVX2 U5 ( .A(s82[3]), .Z(n3) );
  CIVX2 U6 ( .A(c_out800), .Z(n1) );
  CMX2X2 U7 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CND2IX1 U8 ( .B(n1), .A(n5), .Z(n6) );
  CMX2X1 U9 ( .A0(s83[2]), .A1(s84[2]), .S(n8), .Z(sum8[6]) );
  CMX2X2 U10 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CIVXL U11 ( .A(n5), .Z(n4) );
  CMX2XL U12 ( .A0(s83[3]), .A1(s84[3]), .S(n8), .Z(sum8[7]) );
  CMX2X1 U13 ( .A0(s83[1]), .A1(s84[1]), .S(n8), .Z(sum8[5]) );
  CND2XL U14 ( .A(c_in8), .B(c_out801), .Z(n7) );
  CND2X2 U15 ( .A(n6), .B(n7), .Z(n8) );
  CIVXL U16 ( .A(c_in8), .Z(n5) );
  CMX2X2 U17 ( .A0(s83[0]), .A1(s84[0]), .S(n8), .Z(sum8[4]) );
  CMXI2XL U18 ( .A0(n10), .A1(n9), .S(n8), .Z(c_out8) );
  CMXI2X1 U19 ( .A0(n12), .A1(n11), .S(c_in8), .Z(sum8[0]) );
  CIVX2 U20 ( .A(c_out810), .Z(n10) );
  CIVX2 U21 ( .A(c_out811), .Z(n9) );
  CIVX2 U22 ( .A(s81[0]), .Z(n12) );
  CIVX2 U23 ( .A(s82[0]), .Z(n11) );
endmodule


module Add_half_7297 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7298 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3649 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7298 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7297 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7299 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7300 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3650 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7300 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7299 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7301 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7302 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3651 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7302 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7301 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7303 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7304 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3652 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7304 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7303 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_913 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3652 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3651 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3650 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3649 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7305 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7306 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3653 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7306 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7305 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7307 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7308 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3654 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7308 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7307 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7309 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7310 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3655 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7310 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7309 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7311 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7312 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3656 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7312 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7311 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_914 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3656 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3655 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3654 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3653 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7313 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7314 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3657 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7314 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7313 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7315 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7316 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3658 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7316 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7315 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7317 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7318 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3659 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7318 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7317 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7319 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7320 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3660 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7320 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7319 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_915 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3660 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3659 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3658 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3657 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7321 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7322 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3661 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7322 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7321 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7323 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7324 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3662 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7324 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7323 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7325 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7326 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3663 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7326 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7325 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7327 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7328 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3664 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7328 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7327 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_916 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3664 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3663 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3662 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3661 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_229 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_916 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_915 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_914 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_913 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_7329 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7330 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3665 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7330 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7329 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7331 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7332 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3666 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7332 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7331 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7333 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7334 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3667 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7334 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7333 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7335 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7336 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3668 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7336 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7335 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_917 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3668 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3667 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3666 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3665 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7337 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7338 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3669 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7338 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7337 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7339 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7340 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3670 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7340 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7339 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7341 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7342 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3671 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7342 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7341 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7343 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7344 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3672 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7344 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7343 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_918 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3672 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3671 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3670 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3669 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7345 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7346 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3673 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7346 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7345 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7347 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7348 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3674 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7348 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7347 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7349 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7350 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3675 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7350 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7349 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7351 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7352 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3676 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7352 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7351 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_919 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3676 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3675 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3674 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3673 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7353 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7354 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3677 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7354 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7353 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7355 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7356 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3678 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7356 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7355 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7357 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7358 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3679 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7358 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7357 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7359 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7360 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3680 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7360 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7359 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_920 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3680 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3679 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3678 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3677 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_230 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_920 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_919 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_918 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_917 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_7361 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7362 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3681 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7362 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7361 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7363 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7364 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3682 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7364 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7363 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7365 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7366 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3683 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7366 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7365 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7367 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7368 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3684 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7368 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7367 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_921 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3684 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3683 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3682 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3681 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7369 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7370 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3685 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7370 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7369 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7371 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7372 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3686 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7372 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7371 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7373 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7374 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3687 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7374 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7373 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7375 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7376 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3688 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7376 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7375 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_922 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3688 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3687 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3686 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3685 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7377 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7378 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3689 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7378 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7377 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7379 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7380 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3690 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7380 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7379 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7381 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7382 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3691 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7382 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7381 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_7383 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7384 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3692 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7384 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7383 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_923 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_3692 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3691 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3690 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3689 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_7385 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7386 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3693 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7386 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7385 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7387 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7388 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3694 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7388 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7387 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7389 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CENX1 U4 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7390 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3695 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7390 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7389 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7391 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CEOXL U3 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7392 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3696 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7392 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7391 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_924 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_3696 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3695 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3694 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3693 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n4), .A1(n5), .S(n1), .Z(sum2[1]) );
  CMXI2X1 U4 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
endmodule


module bit4_231 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_924 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_923 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_922 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_921 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module Add_half_7393 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7394 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3697 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7394 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7393 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7395 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7396 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3698 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7396 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7395 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7397 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7398 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3699 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7398 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7397 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7399 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7400 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3700 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7400 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7399 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_925 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3700 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3699 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3698 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3697 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7401 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7402 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3701 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7402 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7401 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7403 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7404 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3702 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7404 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7403 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7405 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7406 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3703 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7406 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7405 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7407 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7408 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3704 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7408 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7407 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_926 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3704 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3703 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3702 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3701 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7409 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7410 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3705 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7410 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7409 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7411 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7412 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3706 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7412 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7411 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7413 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7414 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3707 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7414 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7413 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7415 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7416 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3708 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7416 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7415 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_927 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3708 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3707 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3706 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3705 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_7417 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7418 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3709 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7418 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7417 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7419 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7420 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3710 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7420 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7419 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7421 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7422 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3711 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7422 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7421 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7423 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7424 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3712 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7424 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7423 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_928 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3712 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3711 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3710 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3709 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_232 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_928 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_927 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_926 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_925 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CIVX2 U4 ( .A(c_out410), .Z(n3) );
  CIVX2 U5 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n10) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n10), .Z(c_out4) );
  CIVX2 U9 ( .A(s41[0]), .Z(n5) );
  CIVX2 U10 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U12 ( .A(s41[1]), .Z(n7) );
  CIVX2 U13 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U15 ( .A(s43[0]), .Z(n9) );
  CIVX2 U16 ( .A(s44[0]), .Z(n8) );
  CIVX2 U17 ( .A(s43[1]), .Z(n12) );
  CIVX2 U18 ( .A(s44[1]), .Z(n11) );
  CMXI2X1 U19 ( .A0(n12), .A1(n11), .S(n10), .Z(sum4[3]) );
endmodule


module bit8_58 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_232 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_231 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_230 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_229 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CND2X1 U3 ( .A(n6), .B(c_out800), .Z(n7) );
  CND2X1 U4 ( .A(n3), .B(s81[2]), .Z(n4) );
  COR2X1 U5 ( .A(n12), .B(c_in8), .Z(n9) );
  CMX2X1 U6 ( .A0(c_out810), .A1(c_out811), .S(n10), .Z(c_out8) );
  CND2IX1 U7 ( .B(n6), .A(n17), .Z(n18) );
  CANR1XL U8 ( .A(s84[0]), .B(c_out800), .C(n13), .Z(n19) );
  CMXI2X1 U9 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(sum8[1]) );
  CIVX1 U11 ( .A(n6), .Z(n2) );
  CIVX2 U12 ( .A(c_in8), .Z(n6) );
  CMX2X1 U13 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CND2X1 U14 ( .A(c_in8), .B(s82[2]), .Z(n5) );
  CND2X4 U15 ( .A(n4), .B(n5), .Z(sum8[2]) );
  CIVXL U16 ( .A(c_in8), .Z(n3) );
  CND2X1 U17 ( .A(c_in8), .B(c_out801), .Z(n8) );
  CND2X2 U18 ( .A(n7), .B(n8), .Z(n10) );
  CMXI2X1 U19 ( .A0(n23), .A1(n22), .S(n10), .Z(sum8[6]) );
  CMXI2X1 U20 ( .A0(n21), .A1(n20), .S(n10), .Z(sum8[5]) );
  CND2X4 U21 ( .A(n9), .B(n11), .Z(sum8[0]) );
  CND2X1 U22 ( .A(c_in8), .B(s82[0]), .Z(n11) );
  COND1X4 U23 ( .A(n19), .B(n2), .C(n18), .Z(sum8[4]) );
  CNR2IX1 U24 ( .B(s83[0]), .A(c_out800), .Z(n13) );
  CMXI2X2 U25 ( .A0(n25), .A1(n24), .S(n10), .Z(sum8[7]) );
  CIVX2 U26 ( .A(s81[0]), .Z(n12) );
  CIVX2 U27 ( .A(c_out801), .Z(n16) );
  CIVX2 U28 ( .A(s84[0]), .Z(n15) );
  CIVX2 U29 ( .A(s83[0]), .Z(n14) );
  COND2X1 U30 ( .A(n16), .B(n15), .C(c_out801), .D(n14), .Z(n17) );
  CIVX2 U31 ( .A(s83[1]), .Z(n21) );
  CIVX2 U32 ( .A(s84[1]), .Z(n20) );
  CIVX2 U33 ( .A(s83[2]), .Z(n23) );
  CIVX2 U34 ( .A(s84[2]), .Z(n22) );
  CIVX2 U35 ( .A(s83[3]), .Z(n25) );
  CIVX2 U36 ( .A(s84[3]), .Z(n24) );
endmodule


module Add_half_7425 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7426 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3713 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7426 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7425 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7427 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7428 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3714 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7428 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7427 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7429 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7430 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3715 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7430 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7429 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7431 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7432 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3716 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7432 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7431 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_929 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_3716 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3715 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3714 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3713 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_7433 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7434 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3717 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7434 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7433 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7435 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7436 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3718 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7436 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7435 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7437 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7438 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3719 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7438 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7437 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7439 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7440 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3720 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7440 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7439 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_930 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_3720 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3719 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3718 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3717 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_7441 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7442 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3721 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7442 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7441 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7443 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7444 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3722 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7444 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7443 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7445 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7446 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3723 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7446 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7445 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7447 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7448 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3724 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7448 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7447 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_931 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3724 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3723 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3722 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3721 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_7449 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7450 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3725 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7450 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7449 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7451 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7452 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3726 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7452 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7451 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7453 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7454 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3727 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7454 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7453 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7455 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7456 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3728 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7456 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7455 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_932 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3728 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3727 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3726 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3725 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_233 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_932 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_931 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_930 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_929 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2XL U4 ( .A0(n9), .A1(n8), .S(n1), .Z(sum4[3]) );
  CMXI2XL U5 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out4) );
  CMXI2XL U6 ( .A0(n7), .A1(n6), .S(n1), .Z(sum4[2]) );
  CMX2X1 U7 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U8 ( .A(c_out410), .Z(n3) );
  CIVX2 U9 ( .A(c_out411), .Z(n2) );
  CIVX2 U10 ( .A(s41[1]), .Z(n5) );
  CIVX2 U11 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U13 ( .A(s43[0]), .Z(n7) );
  CIVX2 U14 ( .A(s44[0]), .Z(n6) );
  CIVX2 U15 ( .A(s43[1]), .Z(n9) );
  CIVX2 U16 ( .A(s44[1]), .Z(n8) );
endmodule


module Add_half_7457 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7458 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3729 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7458 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7457 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7459 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7460 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3730 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7460 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7459 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7461 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7462 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3731 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7462 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7461 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7463 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7464 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3732 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7464 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7463 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_933 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_3732 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3731 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3730 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3729 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_7465 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7466 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3733 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7466 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7465 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7467 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7468 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3734 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7468 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7467 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7469 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7470 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3735 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7470 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7469 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7471 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7472 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3736 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7472 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7471 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_934 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3736 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3735 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3734 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3733 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVXL U4 ( .A(s3), .Z(n4) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_7473 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7474 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3737 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7474 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7473 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7475 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7476 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3738 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7476 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7475 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7477 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7478 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3739 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7478 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7477 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7479 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7480 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3740 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7480 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7479 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_935 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_3740 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3739 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3738 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3737 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_7481 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7482 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3741 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7482 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7481 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7483 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7484 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3742 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7484 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7483 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7485 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7486 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3743 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7486 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7485 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7487 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7488 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3744 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7488 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7487 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_936 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3744 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3743 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3742 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3741 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_234 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_936 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_935 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_934 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_933 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U7 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
endmodule


module Add_half_7489 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7490 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3745 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7490 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7489 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7491 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7492 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3746 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7492 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7491 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7493 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVXL U1 ( .A(n1), .Z(c_out) );
  CND2XL U2 ( .A(a), .B(b), .Z(n1) );
  CEOXL U3 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7494 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3747 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7494 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7493 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7495 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVXL U1 ( .A(n1), .Z(c_out) );
  CND2XL U2 ( .A(a), .B(b), .Z(n1) );
  CEOXL U3 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7496 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3748 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7496 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7495 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_937 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_3748 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3747 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3746 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3745 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_7497 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CENX1 U4 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7498 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3749 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7498 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7497 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7499 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7500 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3750 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7500 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7499 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7501 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_7502 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3751 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7502 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7501 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7503 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7504 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3752 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7504 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7503 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_938 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3752 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3751 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3750 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3749 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_7505 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CEOXL U3 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7506 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3753 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7506 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7505 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7507 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CEOXL U3 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7508 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3754 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7508 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7507 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7509 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7510 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3755 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7510 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7509 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7511 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7512 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3756 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7512 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7511 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_939 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3756 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3755 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3754 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3753 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_7513 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CENX1 U4 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7514 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3757 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7514 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7513 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7515 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7516 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3758 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7516 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7515 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7517 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7518 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3759 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7518 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7517 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7519 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7520 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3760 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7520 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7519 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_940 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3760 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3759 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3758 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3757 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2XL U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_235 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_940 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_939 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_938 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_937 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module Add_half_7521 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7522 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3761 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7522 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7521 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7523 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7524 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3762 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7524 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7523 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7525 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7526 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3763 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7526 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7525 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7527 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7528 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3764 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7528 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7527 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_941 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3764 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3763 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3762 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3761 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_7529 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_7530 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3765 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7530 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7529 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7531 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7532 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3766 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7532 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7531 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7533 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7534 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3767 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7534 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7533 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7535 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7536 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3768 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7536 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7535 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_942 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3768 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3767 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3766 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3765 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_7537 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7538 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3769 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7538 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7537 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7539 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7540 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3770 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7540 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7539 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7541 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7542 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3771 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7542 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7541 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7543 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7544 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3772 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7544 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7543 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_943 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3772 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3771 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3770 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3769 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_7545 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7546 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3773 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7546 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7545 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7547 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7548 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3774 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7548 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7547 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7549 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7550 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3775 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7550 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7549 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7551 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7552 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3776 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7552 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7551 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_944 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3776 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3775 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3774 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3773 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2XL U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_236 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_944 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_943 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_942 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_941 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CMXI2XL U4 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CMXI2XL U5 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n8) );
  CIVX2 U11 ( .A(s41[1]), .Z(n5) );
  CIVX2 U12 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n7) );
  CIVX2 U15 ( .A(s44[0]), .Z(n6) );
  CIVX2 U16 ( .A(s43[1]), .Z(n10) );
  CIVX2 U17 ( .A(s44[1]), .Z(n9) );
endmodule


module bit8_59 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, net84282, net85320, net85319,
         net90204, net90206, net91091, net93517, n30, net84278, net84810, n1,
         n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;
  assign sum8[0] = net85320;

  bit4_236 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_235 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_234 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_233 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CNR2IX1 U3 ( .B(c_out811), .A(n16), .Z(n1) );
  CIVX2 U4 ( .A(n1), .Z(n7) );
  CND2X1 U5 ( .A(c_out810), .B(n16), .Z(n6) );
  CIVXL U6 ( .A(s84[0]), .Z(n24) );
  CND2X1 U7 ( .A(s81[2]), .B(n2), .Z(n3) );
  CND2XL U8 ( .A(net84810), .B(s82[2]), .Z(n4) );
  CND2X2 U9 ( .A(n3), .B(n4), .Z(sum8[2]) );
  CIVXL U10 ( .A(net84810), .Z(n2) );
  CND2X4 U11 ( .A(n6), .B(n7), .Z(c_out8) );
  CND2X2 U12 ( .A(net84810), .B(s82[0]), .Z(n8) );
  COND1X2 U13 ( .A(net84278), .B(net90206), .C(n8), .Z(n30) );
  CNIVX2 U14 ( .A(c_in8), .Z(net84810) );
  CIVX2 U15 ( .A(net84810), .Z(net84282) );
  CNIVX3 U16 ( .A(c_in8), .Z(net90206) );
  CIVX4 U17 ( .A(n30), .Z(net85319) );
  CIVX2 U18 ( .A(s81[0]), .Z(net84278) );
  CNIVX2 U19 ( .A(net90206), .Z(net90204) );
  CMX2X2 U20 ( .A0(s81[1]), .A1(s82[1]), .S(net90206), .Z(sum8[1]) );
  CND2X4 U21 ( .A(n10), .B(n11), .Z(sum8[6]) );
  CMX2X2 U22 ( .A0(s84[3]), .A1(s83[3]), .S(n14), .Z(sum8[7]) );
  CIVX2 U23 ( .A(n18), .Z(n19) );
  CND2IX2 U24 ( .B(net91091), .A(n23), .Z(n27) );
  CND2X2 U25 ( .A(s84[2]), .B(n9), .Z(n10) );
  CND2X1 U26 ( .A(s83[2]), .B(n15), .Z(n11) );
  CIVX1 U27 ( .A(n15), .Z(n9) );
  COND1X2 U28 ( .A(n25), .B(n20), .C(net90204), .Z(n26) );
  CND2X4 U29 ( .A(n27), .B(n26), .Z(sum8[4]) );
  CND2X2 U30 ( .A(s81[3]), .B(net93517), .Z(n12) );
  CND2X1 U31 ( .A(s82[3]), .B(net90204), .Z(n13) );
  CND2X4 U32 ( .A(n12), .B(n13), .Z(sum8[3]) );
  CIVX1 U33 ( .A(net90204), .Z(net93517) );
  CMXI2X1 U34 ( .A0(n29), .A1(n28), .S(n17), .Z(sum8[5]) );
  CANR2X2 U35 ( .A(net84282), .B(c_out800), .C(n19), .D(net90206), .Z(n16) );
  CANR2XL U36 ( .A(c_out800), .B(net84282), .C(n19), .D(net90206), .Z(n14) );
  CANR2X1 U37 ( .A(net84282), .B(c_out800), .C(n19), .D(net90206), .Z(n15) );
  CANR2X1 U38 ( .A(net84282), .B(c_out800), .C(n19), .D(net90206), .Z(n17) );
  CIVXL U39 ( .A(net84282), .Z(net91091) );
  CIVXL U40 ( .A(c_out801), .Z(n18) );
  CAN2XL U41 ( .A(s84[0]), .B(c_out801), .Z(n20) );
  CIVX8 U42 ( .A(net85319), .Z(net85320) );
  CNR2IXL U43 ( .B(s83[0]), .A(c_out801), .Z(n25) );
  CIVX2 U44 ( .A(c_out800), .Z(n22) );
  CIVX2 U45 ( .A(s83[0]), .Z(n21) );
  COND2X1 U46 ( .A(n22), .B(n24), .C(c_out800), .D(n21), .Z(n23) );
  CIVX2 U47 ( .A(s84[1]), .Z(n29) );
  CIVX2 U48 ( .A(s83[1]), .Z(n28) );
endmodule


module bit32_0 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   n2, c1, c2, c3;

  bit8_0 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8(a32[7:0]), .b8(b32[7:0]), 
        .c_in8(c_in32) );
  bit8_59 A322 ( .sum8(sum32[15:8]), .c_out8(c2), .a8(a32[15:8]), .b8(
        b32[15:8]), .c_in8(c1) );
  bit8_58 A323 ( .sum8({sum32[23:20], n2, sum32[18:16]}), .c_out8(c3), .a8(
        a32[23:16]), .b8(b32[23:16]), .c_in8(c2) );
  bit8_57 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8(a32[31:24]), .b8(
        b32[31:24]), .c_in8(c3) );
  CNIVX4 U1 ( .A(n2), .Z(sum32[19]) );
endmodule


module Add_half_1 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n1) );
  CENX1 U3 ( .A(a), .B(n1), .Z(sum) );
endmodule


module Add_half_2 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_6 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_8 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_4 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_8 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_1 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_4 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0)
         );
  Add_full_3 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1)
         );
  Add_full_2 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0)
         );
  Add_full_1 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1)
         );
  CIVX1 U3 ( .A(n1), .Z(n2) );
  CMX2XL U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_9 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_10 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_5 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_10 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_9 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_11 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_12 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_6 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_12 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_11 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_13 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_14 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_7 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_14 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_13 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_15 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_16 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_8 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_16 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_15 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_2 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n2, n3, n4, n5,
         n6, n7;

  Add_full_8 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0)
         );
  Add_full_7 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1)
         );
  Add_full_6 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0)
         );
  Add_full_5 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1)
         );
  CIVX1 U3 ( .A(s2), .Z(n3) );
  CIVX1 U4 ( .A(s1), .Z(n4) );
  CIVX1 U5 ( .A(s3), .Z(n7) );
  CIVX1 U6 ( .A(s4), .Z(n6) );
  CMXI2X1 U7 ( .A0(n6), .A1(n7), .S(n2), .Z(sum2[1]) );
  CIVDXL U8 ( .A(n2), .Z0(n5) );
  CMX2XL U9 ( .A0(c_out10), .A1(c_out11), .S(n5), .Z(c_out2) );
  CMXI2X1 U10 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMXI2X1 U11 ( .A0(n4), .A1(n3), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_17 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_18 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_9 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_18 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_17 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_19 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_20 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_10 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_20 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_19 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_21 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CNR2X2 U1 ( .A(n1), .B(n2), .Z(c_out) );
  CIVX2 U2 ( .A(a), .Z(n1) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CENXL U4 ( .A(n2), .B(a), .Z(sum) );
endmodule


module Add_half_22 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_11 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_22 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_21 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_23 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CNR2X2 U1 ( .A(n1), .B(n2), .Z(c_out) );
  CIVX2 U2 ( .A(a), .Z(n1) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CEOXL U4 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_24 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4, n5;

  CIVX2 U1 ( .A(b), .Z(n3) );
  CAN2X1 U2 ( .A(b), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(a), .Z(n2) );
  CND2X1 U4 ( .A(a), .B(n3), .Z(n4) );
  CIVXL U5 ( .A(n2), .Z(n1) );
  CND2X2 U6 ( .A(n4), .B(n5), .Z(sum) );
  CND2X2 U7 ( .A(n2), .B(b), .Z(n5) );
endmodule


module Add_full_12 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_24 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_23 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_3 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_12 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_11 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_10 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_9 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1)
         );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX2 U4 ( .A(c_out10), .Z(n4) );
  CIVX2 U5 ( .A(c_out11), .Z(n3) );
  CMX2XL U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U7 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMXI2XL U8 ( .A0(n6), .A1(n5), .S(n1), .Z(sum2[1]) );
  CMX2X1 U9 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module Add_half_25 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_26 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_13 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_26 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_25 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_27 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_28 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_14 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_28 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_27 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_29 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3;

  CNR2X2 U1 ( .A(n1), .B(n2), .Z(c_out) );
  CIVX2 U2 ( .A(a), .Z(n1) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CNIVXL U4 ( .A(a), .Z(n3) );
  CEOXL U5 ( .A(b), .B(n3), .Z(sum) );
endmodule


module Add_half_30 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_15 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_30 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_29 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_31 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3;

  CNIVX1 U1 ( .A(a), .Z(n3) );
  CIVX1 U2 ( .A(a), .Z(n1) );
  CNR2X2 U3 ( .A(n1), .B(n2), .Z(c_out) );
  CIVX2 U4 ( .A(b), .Z(n2) );
  CEOXL U5 ( .A(b), .B(n3), .Z(sum) );
endmodule


module Add_half_32 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X2 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CIVX1 U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_16 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_32 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_31 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_4 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_16 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_15 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_14 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_13 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMX2X2 U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2XL U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U6 ( .A(s2), .Z(n5) );
  CIVX1 U7 ( .A(s1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CIVX2 U9 ( .A(c_out10), .Z(n4) );
  CIVX2 U10 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
endmodule


module bit4_1 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_4 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_3 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_2 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_1 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CND2X1 U3 ( .A(s42[1]), .B(n1), .Z(n2) );
  CND2X2 U4 ( .A(s41[1]), .B(n4), .Z(n3) );
  CND2X2 U5 ( .A(n2), .B(n3), .Z(sum4[1]) );
  CIVX2 U6 ( .A(n4), .Z(n1) );
  CIVX2 U7 ( .A(c_in4), .Z(n4) );
  CIVX2 U8 ( .A(n12), .Z(n5) );
  CND2X2 U9 ( .A(n8), .B(s44[1]), .Z(n9) );
  CIVX2 U10 ( .A(n11), .Z(n8) );
  CND2X2 U11 ( .A(n5), .B(s44[0]), .Z(n6) );
  CND2X1 U12 ( .A(n12), .B(s43[0]), .Z(n7) );
  CND2X2 U13 ( .A(n6), .B(n7), .Z(sum4[2]) );
  CND2X1 U14 ( .A(n11), .B(s43[1]), .Z(n10) );
  CND2X2 U15 ( .A(n9), .B(n10), .Z(sum4[3]) );
  CANR2X1 U16 ( .A(c_out400), .B(n13), .C(c_in4), .D(c_out401), .Z(n11) );
  CANR2X1 U17 ( .A(c_out400), .B(n13), .C(c_in4), .D(c_out401), .Z(n12) );
  CANR2XL U18 ( .A(n13), .B(c_out400), .C(c_in4), .D(c_out401), .Z(n14) );
  CMX2XL U19 ( .A0(c_out411), .A1(c_out410), .S(n14), .Z(c_out4) );
  CMX2X1 U20 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U21 ( .A(c_in4), .Z(n13) );
endmodule


module Add_half_33 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_34 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_17 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_34 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_33 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_35 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n1) );
  CENX1 U3 ( .A(a), .B(n1), .Z(sum) );
endmodule


module Add_half_36 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_18 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_36 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_35 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_37 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(a), .B(n2), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_38 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_19 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_38 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_37 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_39 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(n2) );
  CEOXL U3 ( .A(n2), .B(b), .Z(sum) );
  CAN2X1 U4 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_40 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_20 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_40 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_39 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_5 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_20 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_19 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_18 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_17 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CMX2XL U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CND2X1 U4 ( .A(c_out00), .B(n1), .Z(n2) );
  CND2X1 U5 ( .A(c_out01), .B(c_in2), .Z(n3) );
  CND2X2 U6 ( .A(n2), .B(n3), .Z(n4) );
  CIVX2 U7 ( .A(c_in2), .Z(n1) );
  CMX2XL U8 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMX2X1 U9 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_41 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_42 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_21 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_42 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_41 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_43 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_44 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_22 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_44 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_43 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_45 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_46 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_23 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_46 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_45 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_47 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_48 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_24 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_48 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_47 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_6 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_24 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_23 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_22 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_21 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CDLY1XL U3 ( .A(c_out01), .Z(n1) );
  CMX2X1 U4 ( .A0(c_out00), .A1(n1), .S(c_in2), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CIVXL U6 ( .A(s2), .Z(n4) );
  CIVXL U7 ( .A(s1), .Z(n5) );
  CIVX1 U8 ( .A(s4), .Z(n6) );
  CMXI2X1 U9 ( .A0(n6), .A1(n7), .S(n3), .Z(sum2[1]) );
  CMX2XL U10 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s3), .Z(n7) );
endmodule


module Add_half_49 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_50 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_25 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_50 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_49 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_51 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_52 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_26 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_52 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_51 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_53 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n3;

  CNIVX1 U1 ( .A(a), .Z(n1) );
  CENX1 U2 ( .A(n3), .B(n1), .Z(sum) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U4 ( .A(b), .Z(n3) );
endmodule


module Add_half_54 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_27 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_54 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_53 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_55 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_56 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_28 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_56 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_55 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_7 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11;

  Add_full_28 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_27 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_26 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_25 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CND2X2 U3 ( .A(c_out00), .B(n2), .Z(n3) );
  CMX2X1 U4 ( .A0(n7), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U5 ( .A0(n9), .A1(n8), .S(n5), .Z(c_out2) );
  CND2X2 U6 ( .A(n3), .B(n4), .Z(n5) );
  CIVX1 U7 ( .A(c_out11), .Z(n8) );
  CND2X2 U8 ( .A(c_out01), .B(c_in2), .Z(n4) );
  CIVX2 U9 ( .A(c_in2), .Z(n2) );
  CIVXL U10 ( .A(c_out00), .Z(n6) );
  CIVXL U11 ( .A(n6), .Z(n7) );
  CIVX1 U12 ( .A(c_out10), .Z(n9) );
  CMXI2XL U13 ( .A0(n11), .A1(n10), .S(n1), .Z(sum2[1]) );
  CMX2X1 U14 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U15 ( .A(s3), .Z(n11) );
  CIVX2 U16 ( .A(s4), .Z(n10) );
endmodule


module Add_half_57 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_58 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_29 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_58 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_57 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_59 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_60 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_30 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_60 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_59 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_61 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(n2) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U4 ( .A(b), .B(n2), .Z(sum) );
endmodule


module Add_half_62 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX4 U1 ( .A(b), .Z(n1) );
  CENX2 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_31 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_62 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_61 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_63 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_64 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_32 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_64 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_63 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_8 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_32 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_31 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_30 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_29 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CNIVX1 U3 ( .A(n7), .Z(n1) );
  CIVX2 U4 ( .A(n2), .Z(n7) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX1 U6 ( .A(s2), .Z(n5) );
  CMX2X1 U7 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CIVX1 U8 ( .A(c_out11), .Z(n3) );
  CIVX2 U9 ( .A(c_out10), .Z(n4) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(n7), .Z(c_out2) );
  CIVX2 U11 ( .A(s1), .Z(n6) );
  CMXI2X1 U12 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
endmodule


module bit4_2 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_8 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_7 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_6 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_5 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CND2X1 U3 ( .A(n2), .B(n3), .Z(sum4[2]) );
  CND2X1 U4 ( .A(s44[0]), .B(n1), .Z(n2) );
  CIVX1 U5 ( .A(n7), .Z(n4) );
  CND2X1 U6 ( .A(s43[0]), .B(n8), .Z(n3) );
  CIVX1 U7 ( .A(n8), .Z(n1) );
  CND2X2 U8 ( .A(s44[1]), .B(n4), .Z(n5) );
  CND2X1 U9 ( .A(s43[1]), .B(n7), .Z(n6) );
  CND2X2 U10 ( .A(n6), .B(n5), .Z(sum4[3]) );
  CANR2X1 U11 ( .A(c_out400), .B(n9), .C(c_out401), .D(c_in4), .Z(n7) );
  CANR2X1 U12 ( .A(c_out400), .B(n9), .C(c_in4), .D(c_out401), .Z(n8) );
  CANR2XL U13 ( .A(n9), .B(c_out400), .C(c_in4), .D(c_out401), .Z(n10) );
  CMX2XL U14 ( .A0(c_out411), .A1(c_out410), .S(n10), .Z(c_out4) );
  CMX2X1 U15 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U16 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U17 ( .A(c_in4), .Z(n9) );
endmodule


module Add_half_65 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(n2), .B(a), .Z(sum) );
endmodule


module Add_half_66 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_33 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_66 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_65 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_67 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(n2), .B(a), .Z(sum) );
endmodule


module Add_half_68 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_34 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_68 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_67 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_69 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_70 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_35 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_70 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_69 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_71 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_72 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_36 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_72 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_71 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_9 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_36 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_35 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_34 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_33 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CIVXL U3 ( .A(n1), .Z(n6) );
  CMXI2X1 U4 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_73 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(n2), .B(a), .Z(sum) );
endmodule


module Add_half_74 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_37 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_74 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_73 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_75 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_76 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_38 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_76 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_75 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_77 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_78 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3;

  CND2IX1 U1 ( .B(a), .A(b), .Z(n3) );
  CND2XL U2 ( .A(a), .B(n1), .Z(n2) );
  CND2X1 U3 ( .A(n2), .B(n3), .Z(sum) );
  CIVXL U4 ( .A(b), .Z(n1) );
  CAN2XL U5 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_39 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_78 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_77 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_79 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(n2) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U4 ( .A(b), .B(n2), .Z(sum) );
endmodule


module Add_half_80 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n3), .B(n4), .Z(sum) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n1), .B(b), .Z(n4) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_40 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_80 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_79 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_10 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_40 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_39 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_38 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_37 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CMX2X1 U3 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CIVX2 U4 ( .A(c_in2), .Z(n2) );
  CIVX1 U5 ( .A(c_out10), .Z(n4) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX1 U7 ( .A(s3), .Z(n6) );
  CMXI2XL U8 ( .A0(n6), .A1(n5), .S(n1), .Z(sum2[1]) );
  CIVX2 U9 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(n1), .Z(c_out2) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module Add_half_81 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(a), .B(n2), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_82 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_41 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_82 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_81 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_83 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_84 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_42 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_84 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_83 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_85 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(n1), .Z(sum) );
endmodule


module Add_half_86 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_43 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_86 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_85 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_87 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(n1), .Z(sum) );
endmodule


module Add_half_88 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X2 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X2 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_44 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_88 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_87 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_11 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13;

  Add_full_44 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_43 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_42 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_41 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CMX2X1 U3 ( .A0(n5), .A1(c_out01), .S(c_in2), .Z(n7) );
  CMXI2X1 U4 ( .A0(n13), .A1(n12), .S(n7), .Z(sum2[1]) );
  CMXI2X1 U5 ( .A0(n9), .A1(n8), .S(n3), .Z(c_out2) );
  CND2X2 U6 ( .A(c_out01), .B(c_in2), .Z(n1) );
  CND2X2 U7 ( .A(c_out00), .B(n6), .Z(n2) );
  CND2X2 U8 ( .A(n1), .B(n2), .Z(n3) );
  CIVX2 U9 ( .A(c_in2), .Z(n6) );
  CIVXL U10 ( .A(c_out00), .Z(n4) );
  CIVXL U11 ( .A(n4), .Z(n5) );
  CIVX1 U12 ( .A(s4), .Z(n12) );
  CIVX1 U13 ( .A(s3), .Z(n13) );
  CIVX2 U14 ( .A(c_out10), .Z(n9) );
  CIVX2 U15 ( .A(c_out11), .Z(n8) );
  CIVX2 U16 ( .A(s1), .Z(n11) );
  CIVX2 U17 ( .A(s2), .Z(n10) );
  CMXI2X1 U18 ( .A0(n11), .A1(n10), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_89 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_90 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_45 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_90 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_89 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_91 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CEOXL U3 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_92 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_46 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_92 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_91 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_93 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3;

  CIVXL U1 ( .A(n2), .Z(n1) );
  CNR2X2 U2 ( .A(n2), .B(n3), .Z(c_out) );
  CIVX2 U3 ( .A(a), .Z(n2) );
  CIVX2 U4 ( .A(b), .Z(n3) );
  CENXL U5 ( .A(n3), .B(n1), .Z(sum) );
endmodule


module Add_half_94 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_47 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_94 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_93 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_95 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net85691, n1, n2;
  assign c_out = net85691;

  CNR2X2 U1 ( .A(n1), .B(n2), .Z(net85691) );
  CIVX2 U2 ( .A(a), .Z(n1) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CEOXL U4 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_96 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88016;
  assign c_out = net88016;

  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(net88016) );
endmodule


module Add_full_48 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_96 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_95 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n1), .B(n2), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n2) );
  CIVX2 U3 ( .A(w3), .Z(n1) );
endmodule


module bit2_12 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, net93720,
         net65021, net65020, n1, n2, n3, n4, n5;

  Add_full_48 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_47 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_46 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_45 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CMXI2X1 U3 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CIVX20 U4 ( .A(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n3) );
  CMXI2X1 U6 ( .A0(net65021), .A1(net65020), .S(n2), .Z(c_out2) );
  CIVX2 U7 ( .A(c_out10), .Z(net65020) );
  CIVX2 U8 ( .A(c_out11), .Z(net65021) );
  CMX2XL U9 ( .A0(c_out01), .A1(c_out00), .S(n3), .Z(net93720) );
  CMX2X1 U10 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX1 U11 ( .A(s4), .Z(n4) );
  CIVX1 U12 ( .A(s3), .Z(n5) );
  CMXI2XL U13 ( .A0(n5), .A1(n4), .S(net93720), .Z(sum2[1]) );
endmodule


module bit4_3 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, net65025, net90045, net65033,
         net65032, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_12 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_11 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_10 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_9 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2X1 U4 ( .A0(net65033), .A1(net65032), .S(n1), .Z(c_out4) );
  CMXI2XL U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(net90045) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U7 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX1 U8 ( .A(c_out410), .Z(net65032) );
  CIVX1 U9 ( .A(c_out411), .Z(net65033) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(net65025), .Z(sum4[3]) );
  CIVX1 U11 ( .A(net90045), .Z(net65025) );
  CIVXL U12 ( .A(s43[1]), .Z(n5) );
  CMXI2XL U13 ( .A0(n3), .A1(n2), .S(net65025), .Z(sum4[2]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n3) );
  CIVX2 U15 ( .A(s44[0]), .Z(n2) );
  CIVX2 U16 ( .A(s44[1]), .Z(n4) );
endmodule


module Add_half_97 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_98 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_49 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_98 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_97 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_99 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_100 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_50 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_100 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_99 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_101 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_102 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n1), .B(b), .Z(n4) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CIVXL U3 ( .A(a), .Z(n1) );
  CND2X2 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_51 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_102 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_101 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_103 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U3 ( .A(n1), .B(b), .Z(sum) );
endmodule


module Add_half_104 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_52 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_104 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_103 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_13 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8, n9;

  Add_full_52 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_51 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_50 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_49 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CMXI2XL U3 ( .A0(n9), .A1(n8), .S(n7), .Z(sum2[1]) );
  CIVX1 U4 ( .A(n2), .Z(n7) );
  CIVX2 U5 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CIVX2 U7 ( .A(c_out10), .Z(n4) );
  CIVX2 U8 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n7), .Z(c_out2) );
  CIVX2 U10 ( .A(s1), .Z(n6) );
  CIVX2 U11 ( .A(s2), .Z(n5) );
  CMXI2X1 U12 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U13 ( .A(s3), .Z(n9) );
  CIVX2 U14 ( .A(s4), .Z(n8) );
endmodule


module Add_half_105 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_106 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_53 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_106 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_105 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_107 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_108 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_54 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_108 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_107 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_109 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_110 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_55 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_110 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_109 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_111 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_112 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_56 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_112 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_111 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_14 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_56 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_55 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_54 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_53 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_113 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_114 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(n1), .B(a), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_57 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_114 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_113 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_115 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_116 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_58 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_116 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_115 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_117 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(n2) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U4 ( .A(b), .B(n2), .Z(sum) );
endmodule


module Add_half_118 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX2 U1 ( .A(n1), .B(a), .Z(sum) );
  CIVX4 U2 ( .A(b), .Z(n1) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_59 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_118 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_117 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_119 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CNR2X2 U1 ( .A(n1), .B(n2), .Z(c_out) );
  CIVX2 U2 ( .A(a), .Z(n1) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CEOXL U4 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_120 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_60 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_120 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_119 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_15 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8, n9;

  Add_full_60 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_59 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_58 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_57 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CIVX2 U4 ( .A(c_out11), .Z(n4) );
  CMXI2X1 U5 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n3) );
  CIVX1 U6 ( .A(s4), .Z(n8) );
  CIVX1 U7 ( .A(s3), .Z(n9) );
  CIVX1 U8 ( .A(s2), .Z(n6) );
  CIVX1 U9 ( .A(s1), .Z(n7) );
  CMX2XL U10 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMXI2X1 U11 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CIVX2 U12 ( .A(c_out10), .Z(n5) );
  CMXI2X1 U13 ( .A0(n7), .A1(n6), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U14 ( .A0(n9), .A1(n8), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_121 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_122 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_61 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_122 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_121 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_123 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_124 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_62 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_124 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_123 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_125 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(a), .B(n2), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_126 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVXL U1 ( .A(b), .Z(n2) );
  CND2X1 U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CND2X1 U4 ( .A(n1), .B(b), .Z(n4) );
  CIVX1 U5 ( .A(a), .Z(n1) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_63 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_126 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_125 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_127 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_128 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X2 U1 ( .A(n1), .B(b), .Z(n4) );
  CIVX2 U2 ( .A(a), .Z(n1) );
  CND2X1 U3 ( .A(a), .B(n2), .Z(n3) );
  CND2X2 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_64 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_128 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_127 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_16 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_64 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_63 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_62 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_61 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CND2X2 U3 ( .A(c_out01), .B(c_in2), .Z(n3) );
  CMXI2X1 U4 ( .A0(n7), .A1(n6), .S(n4), .Z(c_out2) );
  CND2X2 U5 ( .A(c_out00), .B(n1), .Z(n2) );
  CND2X2 U6 ( .A(n2), .B(n3), .Z(n4) );
  CIVX2 U7 ( .A(c_in2), .Z(n1) );
  CMX2XL U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n5) );
  CIVX1 U9 ( .A(c_out10), .Z(n7) );
  CMX2XL U10 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U11 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(c_out11), .Z(n6) );
endmodule


module bit4_4 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_16 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_15 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_14 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_13 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(c_out411), .Z(n4) );
  CMX2X2 U4 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CIVX2 U5 ( .A(c_in4), .Z(n1) );
  CMX2X1 U6 ( .A0(s43[0]), .A1(s44[0]), .S(n2), .Z(sum4[2]) );
  CMXI2X1 U7 ( .A0(c_out401), .A1(c_out400), .S(n1), .Z(n3) );
  CIVX1 U8 ( .A(c_out410), .Z(n5) );
  CMXI2X1 U9 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out4) );
  CMX2X1 U10 ( .A0(s43[1]), .A1(s44[1]), .S(n2), .Z(sum4[3]) );
  CMX2X1 U11 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U12 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
endmodule


module bit8_1 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, net65177, net89993, net90429,
         net93174, net93253, net65176, net65175, net65179, net65178, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_4 A81 ( .sum4(s81), .c_out4(c_out800), .a4({a8[3:1], n5}), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_3 A82 ( .sum4(s82), .c_out4(c_out801), .a4({a8[3:1], n6}), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_2 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4({b8[7:5], n8}), 
        .c_in4(1'b0) );
  bit4_1 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4({b8[7:5], n8}), 
        .c_in4(1'b1) );
  CIVX1 U3 ( .A(s83[2]), .Z(net65179) );
  CIVX1 U4 ( .A(n3), .Z(net90429) );
  CIVX2 U5 ( .A(n2), .Z(n1) );
  CIVXL U6 ( .A(net93253), .Z(n2) );
  CIVX1 U7 ( .A(s81[2]), .Z(n12) );
  CMXI2X1 U8 ( .A0(n11), .A1(n12), .S(net93253), .Z(sum8[2]) );
  CMX2X1 U9 ( .A0(s81[3]), .A1(s82[3]), .S(net90429), .Z(sum8[3]) );
  CIVX1 U10 ( .A(net90429), .Z(net93253) );
  CMX2X1 U11 ( .A0(s82[1]), .A1(s81[1]), .S(net93174), .Z(sum8[1]) );
  CMXI2X1 U12 ( .A0(net65178), .A1(net65179), .S(n4), .Z(sum8[6]) );
  CIVX2 U13 ( .A(s84[2]), .Z(net65178) );
  CANR2X1 U14 ( .A(n3), .B(c_out800), .C(c_in8), .D(c_out801), .Z(n4) );
  CMXI2X1 U15 ( .A0(net65175), .A1(net65176), .S(n4), .Z(sum8[7]) );
  CIVX2 U16 ( .A(c_in8), .Z(n3) );
  CANR2X1 U17 ( .A(n3), .B(c_out800), .C(c_in8), .D(c_out801), .Z(net65177) );
  CANR2XL U18 ( .A(n1), .B(c_out800), .C(n2), .D(c_out801), .Z(net89993) );
  CIVXL U19 ( .A(c_in8), .Z(net93174) );
  CNIVX4 U20 ( .A(a8[0]), .Z(n5) );
  CNIVX4 U21 ( .A(a8[0]), .Z(n6) );
  CIVX2 U22 ( .A(s83[3]), .Z(net65176) );
  CIVX2 U23 ( .A(s84[3]), .Z(net65175) );
  CMX2X1 U24 ( .A0(s81[0]), .A1(s82[0]), .S(net90429), .Z(sum8[0]) );
  CIVXL U25 ( .A(s82[2]), .Z(n11) );
  CIVX8 U26 ( .A(n7), .Z(n8) );
  CIVX2 U27 ( .A(b8[4]), .Z(n7) );
  CMXI2XL U28 ( .A0(n10), .A1(n9), .S(net89993), .Z(c_out8) );
  CIVX2 U29 ( .A(c_out811), .Z(n10) );
  CIVX2 U30 ( .A(c_out810), .Z(n9) );
  CIVX2 U31 ( .A(s84[0]), .Z(n14) );
  CIVX2 U32 ( .A(s83[0]), .Z(n13) );
  CMXI2X1 U33 ( .A0(n14), .A1(n13), .S(net65177), .Z(sum8[4]) );
  CIVX2 U34 ( .A(s84[1]), .Z(n16) );
  CIVX2 U35 ( .A(s83[1]), .Z(n15) );
  CMXI2X1 U36 ( .A0(n16), .A1(n15), .S(net65177), .Z(sum8[5]) );
endmodule


module Add_half_129 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_130 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_65 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_130 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_129 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_131 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_132 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_66 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_132 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_131 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_133 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CEOXL U3 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_134 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_67 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_134 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_133 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_135 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_136 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_68 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_136 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_135 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_17 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_68 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_67 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_66 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_65 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_137 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_138 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_69 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_138 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_137 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_139 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_140 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_70 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_140 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_139 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_141 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_142 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_71 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_142 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_141 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_143 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_144 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVX1 U1 ( .A(a), .Z(n1) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_72 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_144 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_143 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_18 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_72 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_71 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_70 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_69 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n3), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n3), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(n2), .Z(n3) );
endmodule


module Add_half_145 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_146 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_73 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_146 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_145 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_147 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_148 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_74 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_148 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_147 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_149 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CDLY1X2 U1 ( .A(a), .Z(n1) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(n1), .Z(sum) );
endmodule


module Add_half_150 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_75 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_150 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_149 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_151 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X2 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_152 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_76 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_152 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_151 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X2 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_19 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10;

  Add_full_76 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_75 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_74 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_73 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CMXI2X1 U3 ( .A0(n10), .A1(n9), .S(n2), .Z(sum2[1]) );
  CDLY1XL U4 ( .A(c_out01), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n3) );
  CMX2XL U6 ( .A0(n1), .A1(c_out00), .S(n3), .Z(n2) );
  CMXI2X1 U7 ( .A0(n5), .A1(n6), .S(n4), .Z(c_out2) );
  CMXI2X1 U8 ( .A0(c_out01), .A1(c_out00), .S(n3), .Z(n4) );
  CIVX2 U9 ( .A(c_out10), .Z(n6) );
  CIVX2 U10 ( .A(c_out11), .Z(n5) );
  CIVX2 U11 ( .A(s1), .Z(n8) );
  CIVX2 U12 ( .A(s2), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U14 ( .A(s3), .Z(n10) );
  CIVX2 U15 ( .A(s4), .Z(n9) );
endmodule


module Add_half_153 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(a), .B(n2), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_154 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_77 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_154 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_153 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_155 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_156 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_78 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_156 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_155 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_157 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_158 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_79 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_158 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_157 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_159 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CDLY1XL U2 ( .A(a), .Z(n2) );
  CEOXL U3 ( .A(n2), .B(b), .Z(sum) );
endmodule


module Add_half_160 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_80 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_160 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_159 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_20 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_80 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_79 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_78 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_77 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out10), .Z(n4) );
  CIVX2 U9 ( .A(c_out11), .Z(n3) );
endmodule


module bit4_5 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_20 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_19 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_18 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_17 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(n5), .Z(n8) );
  CMXI2X1 U4 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n5) );
  CND2X2 U5 ( .A(n3), .B(n4), .Z(c_out4) );
  CND2X1 U6 ( .A(n8), .B(c_out411), .Z(n4) );
  CIVXL U7 ( .A(n2), .Z(n1) );
  CIVX2 U8 ( .A(n8), .Z(n2) );
  CND2X2 U9 ( .A(c_out410), .B(n2), .Z(n3) );
  CMX2XL U10 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U11 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U12 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMXI2XL U13 ( .A0(n7), .A1(n6), .S(n1), .Z(sum4[2]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n7) );
  CIVX2 U15 ( .A(s44[0]), .Z(n6) );
endmodule


module Add_half_161 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_162 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_81 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_162 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_161 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_163 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_164 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_82 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_164 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_163 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_165 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_166 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_83 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_166 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_165 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_167 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_168 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_84 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_168 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_167 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_21 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_84 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_83 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_82 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_81 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CIVX1 U4 ( .A(n2), .Z(n5) );
  CMXI2X1 U5 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(c_out10), .A1(c_out11), .S(n5), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n4) );
  CIVX2 U9 ( .A(s2), .Z(n3) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_169 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_170 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_85 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_170 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_169 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_171 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_172 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_86 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_172 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_171 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_173 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_174 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_87 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_174 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_173 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_175 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_176 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_88 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_176 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_175 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_22 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_88 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_87 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_86 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_85 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CMXI2X1 U3 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n3) );
  CIVX20 U4 ( .A(c_in2), .Z(n1) );
  CMX2XL U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMX2X1 U6 ( .A0(c_out11), .A1(c_out10), .S(n3), .Z(c_out2) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(s3), .Z(n5) );
  CIVX2 U9 ( .A(s4), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_177 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_178 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_89 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_178 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_177 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_179 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_180 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_90 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_180 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_179 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_181 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CDLY1X2 U3 ( .A(a), .Z(n2) );
  CEOXL U4 ( .A(b), .B(n2), .Z(sum) );
endmodule


module Add_half_182 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_91 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_182 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_181 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_183 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CDLY1XL U1 ( .A(a), .Z(n1) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(n1), .Z(sum) );
endmodule


module Add_half_184 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_92 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_184 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_183 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_23 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_92 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_91 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_90 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_89 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CIVX1 U4 ( .A(c_out10), .Z(n5) );
  CIVX1 U5 ( .A(c_out11), .Z(n4) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n3) );
  CIVX1 U7 ( .A(s1), .Z(n7) );
  CMX2XL U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMXI2X1 U9 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CMX2XL U10 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CIVX2 U11 ( .A(s2), .Z(n6) );
  CMXI2X1 U12 ( .A0(n7), .A1(n6), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_185 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_186 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_93 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_186 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_185 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_187 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_188 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_94 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_188 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_187 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_189 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n3;

  CENX1 U1 ( .A(n3), .B(n1), .Z(sum) );
  CDLY1XL U2 ( .A(a), .Z(n1) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U4 ( .A(b), .Z(n3) );
endmodule


module Add_half_190 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_95 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_190 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_189 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_191 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CDLY1XL U1 ( .A(a), .Z(n1) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(n1), .Z(sum) );
endmodule


module Add_half_192 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_96 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_192 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_191 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_24 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8, n9;

  Add_full_96 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(1'b0) );
  Add_full_95 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_94 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_93 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CIVXL U3 ( .A(c_out00), .Z(n1) );
  CIVXL U4 ( .A(n1), .Z(n2) );
  CMX2XL U5 ( .A0(n2), .A1(c_out01), .S(c_in2), .Z(n3) );
  CIVX2 U6 ( .A(c_in2), .Z(n4) );
  CMXI2X1 U7 ( .A0(c_out01), .A1(c_out00), .S(n4), .Z(n5) );
  CMXI2X1 U8 ( .A0(n6), .A1(n7), .S(n5), .Z(c_out2) );
  CMX2X1 U9 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2XL U10 ( .A0(n9), .A1(n8), .S(n3), .Z(sum2[1]) );
  CIVX2 U11 ( .A(c_out10), .Z(n7) );
  CIVX2 U12 ( .A(c_out11), .Z(n6) );
  CIVX2 U13 ( .A(s3), .Z(n9) );
  CIVX2 U14 ( .A(s4), .Z(n8) );
endmodule


module bit4_6 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_24 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_23 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_22 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_21 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVXL U3 ( .A(n6), .Z(n2) );
  CIVX1 U4 ( .A(c_out411), .Z(n7) );
  CIVX2 U5 ( .A(n2), .Z(n1) );
  CIVX1 U6 ( .A(c_out410), .Z(n8) );
  CND2X1 U7 ( .A(c_out400), .B(n3), .Z(n4) );
  CND2X1 U8 ( .A(c_out401), .B(c_in4), .Z(n5) );
  CND2X2 U9 ( .A(n4), .B(n5), .Z(n6) );
  CIVX2 U10 ( .A(c_in4), .Z(n3) );
  CMX2XL U11 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2XL U12 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2X1 U13 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U14 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMXI2X1 U15 ( .A0(n8), .A1(n7), .S(n6), .Z(c_out4) );
endmodule


module Add_half_193 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CEOXL U3 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_194 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_97 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_194 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_193 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_195 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CENX1 U4 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_196 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_98 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_196 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_195 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_197 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_198 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_99 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_198 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_197 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_199 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_200 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net89368;
  assign c_out = net89368;

  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(net89368) );
endmodule


module Add_full_100 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_200 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_199 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_25 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, net65502,
         net65503, net65501, n1, n2, n3, n4;

  Add_full_100 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_99 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(1'b1) );
  Add_full_98 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(1'b0) );
  Add_full_97 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(1'b1) );
  CIVX1 U3 ( .A(n3), .Z(net65501) );
  CIVX2 U4 ( .A(c_in2), .Z(n4) );
  CMXI2X1 U5 ( .A0(n1), .A1(n2), .S(net65501), .Z(c_out2) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n4), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CIVX2 U8 ( .A(c_out10), .Z(n1) );
  CMXI2X1 U9 ( .A0(net65502), .A1(net65503), .S(c_in2), .Z(sum2[0]) );
  CMX2XL U10 ( .A0(s3), .A1(s4), .S(net65501), .Z(sum2[1]) );
  CIVX2 U11 ( .A(s1), .Z(net65502) );
  CIVX2 U12 ( .A(s2), .Z(net65503) );
endmodule


module Add_half_201 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_202 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_101 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_202 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_201 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_203 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_204 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_102 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_204 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_203 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_205 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n3;

  CDLY1XL U1 ( .A(a), .Z(n1) );
  CENXL U2 ( .A(n1), .B(n3), .Z(sum) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U4 ( .A(b), .Z(n3) );
endmodule


module Add_half_206 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3;

  CIVX1 U1 ( .A(a), .Z(n1) );
  CND2X1 U2 ( .A(n3), .B(n2), .Z(sum) );
  CND2IXL U3 ( .B(b), .A(a), .Z(n2) );
  CND2X1 U4 ( .A(n1), .B(b), .Z(n3) );
  CAN2XL U5 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_103 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_206 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_205 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_207 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CDLY1XL U1 ( .A(a), .Z(n1) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(n1), .Z(sum) );
endmodule


module Add_half_208 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_104 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_208 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_207 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_26 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_104 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_103 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_102 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_101 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CNIVXL U3 ( .A(n3), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMXI2XL U5 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CIVX1 U6 ( .A(n2), .Z(n3) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMX2X1 U8 ( .A0(c_out10), .A1(c_out11), .S(n3), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
endmodule


module Add_half_209 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_210 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_105 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_210 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_209 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_211 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_212 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_106 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_212 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_211 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_213 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_214 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X2 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X2 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX2 U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_107 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_214 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_213 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_215 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n3;

  CND2IX2 U1 ( .B(n3), .A(a), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CENXL U3 ( .A(n3), .B(a), .Z(sum) );
  CIVX2 U4 ( .A(b), .Z(n3) );
endmodule


module Add_half_216 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88836, n1, n2, n3, n4;
  assign c_out = net88836;

  CIVX1 U1 ( .A(a), .Z(n1) );
  CND2XL U2 ( .A(n2), .B(a), .Z(n3) );
  CND2X2 U3 ( .A(n1), .B(b), .Z(n4) );
  CND2X2 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(net88836) );
endmodule


module Add_full_108 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_216 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_215 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_27 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, net95635,
         net65569, net65568, n1;

  Add_full_108 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_107 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_106 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_105 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(net65569), .A1(net65568), .S(n1), .Z(c_out2) );
  CMXI2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(c_out10), .Z(net65568) );
  CIVX2 U6 ( .A(c_out11), .Z(net65569) );
  CMX2XL U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(net95635) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMX2XL U9 ( .A0(s3), .A1(s4), .S(net95635), .Z(sum2[1]) );
endmodule


module Add_half_217 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_218 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_109 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_218 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_217 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_219 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_220 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_110 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_220 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_219 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_221 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net86446, n1, n2, n3;
  assign c_out = net86446;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CEOXL U2 ( .A(n3), .B(b), .Z(sum) );
  CND2IX1 U3 ( .B(n1), .A(a), .Z(n2) );
  CNIVXL U4 ( .A(a), .Z(n3) );
  CIVX2 U5 ( .A(n2), .Z(net86446) );
endmodule


module Add_half_222 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88833;
  assign c_out = net88833;

  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(net88833) );
endmodule


module Add_full_111 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_222 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_221 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_223 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net86447, n1, n2, n3;
  assign c_out = net86447;

  CND2IX1 U1 ( .B(n1), .A(a), .Z(n2) );
  CIVX2 U2 ( .A(b), .Z(n1) );
  CIVX2 U3 ( .A(n2), .Z(net86447) );
  CDLY1X2 U4 ( .A(a), .Z(n3) );
  CEOX2 U5 ( .A(n3), .B(b), .Z(sum) );
endmodule


module Add_half_224 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88834;
  assign c_out = net88834;

  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(net88834) );
endmodule


module Add_full_112 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_224 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_223 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_28 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, net65598,
         net65599, net95755, net65597, n1, n2, n3, n4, n5;

  Add_full_112 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_111 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_110 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_109 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n5), .A1(n4), .S(net95755), .Z(sum2[1]) );
  CMXI2X1 U4 ( .A0(n1), .A1(n2), .S(net65597), .Z(c_out2) );
  CIVX2 U5 ( .A(n3), .Z(net65597) );
  CDLY1XL U6 ( .A(net65597), .Z(net95755) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CIVX2 U9 ( .A(c_out10), .Z(n1) );
  CMXI2X1 U10 ( .A0(net65598), .A1(net65599), .S(c_in2), .Z(sum2[0]) );
  CIVX1 U11 ( .A(s2), .Z(net65599) );
  CIVX1 U12 ( .A(s1), .Z(net65598) );
  CIVX2 U13 ( .A(s3), .Z(n5) );
  CIVX2 U14 ( .A(s4), .Z(n4) );
endmodule


module bit4_7 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, net100822, net65613, net65612,
         n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_28 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_27 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_26 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_25 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVXL U3 ( .A(c_out400), .Z(n1) );
  CIVXL U4 ( .A(n1), .Z(n2) );
  CIVXL U5 ( .A(c_out401), .Z(n3) );
  CIVXL U6 ( .A(n3), .Z(n4) );
  CIVX2 U7 ( .A(c_in4), .Z(n5) );
  CMXI2X1 U8 ( .A0(c_out401), .A1(c_out400), .S(n5), .Z(n6) );
  CMXI2X1 U9 ( .A0(net65613), .A1(net65612), .S(n6), .Z(c_out4) );
  CMX2XL U10 ( .A0(n2), .A1(n4), .S(c_in4), .Z(net100822) );
  CMX2X1 U11 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U12 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX1 U13 ( .A(c_out410), .Z(net65612) );
  CIVX1 U14 ( .A(c_out411), .Z(net65613) );
  CMX2XL U15 ( .A0(s43[1]), .A1(s44[1]), .S(net100822), .Z(sum4[3]) );
  CMX2XL U16 ( .A0(s43[0]), .A1(s44[0]), .S(net100822), .Z(sum4[2]) );
endmodule


module Add_half_225 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CEOXL U3 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_226 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_113 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_226 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_225 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_227 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CEOXL U3 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_228 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_114 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_228 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_227 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_229 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_230 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_115 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_230 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_229 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_231 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_232 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(a), .B(n2), .Z(n3) );
  CIVX1 U2 ( .A(a), .Z(n1) );
  CND2X1 U3 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_116 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_232 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_231 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_29 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_116 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_115 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_114 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_113 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s3), .Z(n8) );
  CIVX2 U13 ( .A(s4), .Z(n7) );
endmodule


module Add_half_233 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CENX1 U4 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_234 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_117 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_234 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_233 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_235 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_236 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_118 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_236 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_235 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_237 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_238 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_119 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_238 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_237 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_239 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_240 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(a), .B(n2), .Z(n3) );
  CIVX1 U2 ( .A(a), .Z(n1) );
  CND2X1 U3 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_120 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_240 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_239 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_30 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_120 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_119 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_118 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_117 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_241 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_242 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_121 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_242 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_241 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_243 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_244 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_122 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_244 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_243 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_245 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_246 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_123 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_246 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_245 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_247 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_248 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_124 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_248 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_247 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_31 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10;

  Add_full_124 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_123 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_122 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_121 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(n8), .Z(n1) );
  CIVXL U4 ( .A(n1), .Z(n2) );
  CIVX1 U5 ( .A(s2), .Z(n6) );
  CMXI2XL U6 ( .A0(n10), .A1(n9), .S(n2), .Z(sum2[1]) );
  CIVX2 U7 ( .A(n3), .Z(n8) );
  CIVX1 U8 ( .A(s1), .Z(n7) );
  CIVX2 U9 ( .A(c_out10), .Z(n5) );
  CIVX2 U10 ( .A(c_out11), .Z(n4) );
  CMXI2X1 U11 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(n8), .Z(c_out2) );
  CMXI2X1 U13 ( .A0(n7), .A1(n6), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U14 ( .A(s3), .Z(n10) );
  CIVX2 U15 ( .A(s4), .Z(n9) );
endmodule


module Add_half_249 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_250 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_125 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_250 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_249 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_251 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_252 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_126 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_252 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_251 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_253 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_254 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_127 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_254 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_253 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_255 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_256 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_full_128 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_256 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_255 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_32 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_128 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_127 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_126 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_125 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_8 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_32 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_31 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_30 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_29 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out4) );
  CIVXL U4 ( .A(n1), .Z(n4) );
  CIVX1 U5 ( .A(c_out411), .Z(n2) );
  CIVX1 U6 ( .A(c_out410), .Z(n3) );
  CMX2XL U7 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2XL U8 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U9 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U10 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMXI2X1 U11 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
endmodule


module bit8_2 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, net90004, net90003, net90268,
         net90267, net90277, net90276, net91184, net91182, n1, n2, n3, n4, n5,
         n6, n7, n8;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_8 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_7 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_6 A83 ( .sum4(s83), .c_out4(c_out810), .a4({a8[7:5], n7}), .b4({n8, 
        b8[6:5], n4}), .c_in4(1'b0) );
  bit4_5 A84 ( .sum4(s84), .c_out4(c_out811), .a4({a8[7:5], n5}), .b4({n8, 
        b8[6:5], n4}), .c_in4(1'b1) );
  CIVX2 U3 ( .A(n6), .Z(n5) );
  CIVX1 U4 ( .A(a8[4]), .Z(n6) );
  CIVX2 U5 ( .A(c_in8), .Z(n2) );
  CND2X2 U6 ( .A(n3), .B(net91184), .Z(c_out8) );
  CND2X1 U7 ( .A(n1), .B(c_out810), .Z(net91184) );
  CND2X2 U8 ( .A(net91182), .B(c_out811), .Z(n3) );
  CIVX2 U9 ( .A(n1), .Z(net91182) );
  CANR2X2 U10 ( .A(n2), .B(c_out800), .C(c_in8), .D(c_out801), .Z(n1) );
  CANR2XL U11 ( .A(net90277), .B(n2), .C(c_in8), .D(net90268), .Z(net90004) );
  CANR2XL U12 ( .A(n2), .B(net90277), .C(c_in8), .D(net90268), .Z(net90003) );
  CIVXL U13 ( .A(c_out800), .Z(net90276) );
  CIVXL U14 ( .A(c_out801), .Z(net90267) );
  CNIVX4 U15 ( .A(b8[4]), .Z(n4) );
  CIVX1 U16 ( .A(n6), .Z(n7) );
  CIVXL U17 ( .A(net90276), .Z(net90277) );
  CIVXL U18 ( .A(net90267), .Z(net90268) );
  CNIVX4 U19 ( .A(b8[7]), .Z(n8) );
  CMX2XL U20 ( .A0(s84[2]), .A1(s83[2]), .S(net90004), .Z(sum8[6]) );
  CMX2XL U21 ( .A0(s84[3]), .A1(s83[3]), .S(net90003), .Z(sum8[7]) );
  CMX2XL U22 ( .A0(s84[0]), .A1(s83[0]), .S(net90004), .Z(sum8[4]) );
  CMX2XL U23 ( .A0(s84[1]), .A1(s83[1]), .S(net90003), .Z(sum8[5]) );
  CMX2XL U24 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2XL U25 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2XL U26 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2XL U27 ( .A0(s81[0]), .A1(s82[0]), .S(c_in8), .Z(sum8[0]) );
endmodule


module Add_half_257 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_258 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_129 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_258 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_257 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_259 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_260 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_130 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_260 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_259 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_261 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_262 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_131 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_262 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_261 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_263 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_264 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_132 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_264 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_263 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_33 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_132 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_131 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_130 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_129 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_265 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_266 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_133 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_266 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_265 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_267 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_268 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_134 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_268 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_267 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_269 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_270 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_135 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_270 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_269 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_271 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_272 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_136 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_272 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_271 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_34 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_136 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_135 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_134 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_133 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module Add_half_273 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_274 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_137 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_274 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_273 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_275 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_276 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_138 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_276 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_275 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_277 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_278 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_139 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_278 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_277 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_279 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_280 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_140 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_280 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_279 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_35 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n2, n3, n4, n5,
         n6, n7, n8, n9;

  Add_full_140 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_139 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_138 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_137 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CIVDXL U4 ( .A(n2), .Z0(n7) );
  CIVX2 U5 ( .A(c_out10), .Z(n4) );
  CIVX2 U6 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX2 U8 ( .A(s1), .Z(n6) );
  CIVX2 U9 ( .A(s2), .Z(n5) );
  CMXI2X1 U10 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n9) );
  CIVX2 U12 ( .A(s4), .Z(n8) );
  CMXI2X1 U13 ( .A0(n9), .A1(n8), .S(n7), .Z(sum2[1]) );
endmodule


module Add_half_281 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_282 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_141 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_282 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_281 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_283 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_284 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_142 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_284 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_283 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_285 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_286 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_143 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_286 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_285 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_287 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_288 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_144 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_288 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_287 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_36 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_144 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_143 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_142 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_141 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_9 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_36 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_35 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_34 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_33 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CND2XL U3 ( .A(c_out410), .B(n1), .Z(n2) );
  CND2XL U4 ( .A(c_out411), .B(n4), .Z(n3) );
  CND2X1 U5 ( .A(n2), .B(n3), .Z(c_out4) );
  CIVXL U6 ( .A(n4), .Z(n1) );
  CMX2XL U7 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n4) );
  CMX2XL U9 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U10 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U11 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
endmodule


module Add_half_289 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_290 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_145 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_290 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_289 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_291 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_292 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_146 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_292 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_291 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_293 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVX1 U1 ( .A(a), .Z(n1) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(n1), .Z(sum) );
endmodule


module Add_half_294 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_147 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_294 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_293 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_295 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_296 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_148 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_296 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_295 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_37 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_148 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_147 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_146 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_145 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s1), .Z(n3) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CIVX2 U7 ( .A(s2), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_297 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_298 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_149 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_298 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_297 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_299 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_300 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_150 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_300 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_299 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_301 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_302 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_151 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_302 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_301 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_303 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_304 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_152 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_304 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_303 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_38 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_152 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_151 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_150 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_149 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_305 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_306 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_153 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_306 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_305 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_307 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_308 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_154 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_308 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_307 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_309 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_310 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_155 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_310 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_309 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_311 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_312 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_156 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_312 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_311 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_39 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_156 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_155 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_154 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_153 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2XL U4 ( .A0(n7), .A1(n6), .S(n1), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n7) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
endmodule


module Add_half_313 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_314 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_157 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_314 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_313 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_315 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_316 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_158 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_316 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_315 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_317 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_318 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_159 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_318 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_317 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_319 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_320 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_160 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_320 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_319 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_40 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_160 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_159 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_158 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_157 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n4) );
  CIVX2 U8 ( .A(c_out11), .Z(n3) );
  CIVX2 U9 ( .A(n2), .Z(n5) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(n5), .Z(c_out2) );
endmodule


module bit4_10 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_40 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_39 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_38 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_37 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX1 U7 ( .A(c_out411), .Z(n2) );
  CIVX1 U8 ( .A(c_out410), .Z(n3) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module Add_half_321 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_322 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_161 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_322 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_321 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_323 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_324 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_162 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_324 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_323 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_325 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_326 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_163 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_326 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_325 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_327 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_328 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVXL U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_164 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_328 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_327 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_41 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_164 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_163 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_162 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_161 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMXI2X1 U3 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CMXI2XL U4 ( .A0(n4), .A1(n5), .S(n1), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module Add_half_329 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_330 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_165 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_330 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_329 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_331 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_332 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_166 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_332 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_331 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_333 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_334 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_167 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_334 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_333 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_335 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_336 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_168 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_336 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_335 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_42 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_168 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_167 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_166 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_165 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CMXI2XL U3 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX1 U4 ( .A(n1), .Z(n4) );
  CIVX1 U5 ( .A(s3), .Z(n6) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_337 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_338 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_169 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_338 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_337 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_339 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_340 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_170 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_340 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_339 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_341 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_342 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_171 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_342 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_341 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_343 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(n2) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U4 ( .A(b), .B(n2), .Z(sum) );
endmodule


module Add_half_344 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_172 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_344 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_343 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_43 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_172 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_171 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_170 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_169 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_345 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_346 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_173 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_346 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_345 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_347 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_348 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_174 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_348 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_347 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_349 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_350 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_175 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_350 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_349 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_351 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_352 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_176 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_352 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_351 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_44 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_176 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_175 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_174 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_173 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CIVX1 U4 ( .A(s3), .Z(n6) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module bit4_11 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_44 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_43 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_42 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_41 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CIVX1 U3 ( .A(c_out411), .Z(n2) );
  CIVX1 U4 ( .A(c_out410), .Z(n3) );
  CMX2XL U5 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2XL U6 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2X1 U7 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMX2X1 U8 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out4) );
  CIVX2 U11 ( .A(c_in4), .Z(n4) );
endmodule


module Add_half_353 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_354 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_177 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_354 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_353 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_355 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_356 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_178 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_356 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_355 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_357 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_358 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_179 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_358 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_357 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_359 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_360 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_180 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_360 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_359 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_45 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_180 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_179 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_178 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_177 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CMXI2XL U3 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX1 U4 ( .A(n1), .Z(n4) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_361 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_362 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_181 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_362 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_361 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_363 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_364 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_182 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_364 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_363 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_365 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_366 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_183 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_366 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_365 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_367 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_368 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_184 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_368 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_367 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_46 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_184 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_183 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_182 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_181 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVXL U3 ( .A(s3), .Z(n6) );
  CMXI2XL U4 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n4) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_369 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_370 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_185 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_370 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_369 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_371 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_372 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_186 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_372 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_371 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_373 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_374 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_187 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_374 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_373 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_375 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_376 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_188 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_376 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_375 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_47 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_188 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_187 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_186 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_185 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_377 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_378 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_189 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_378 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_377 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_379 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_380 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_190 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_380 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_379 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_381 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_382 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_191 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_382 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_381 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_383 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_384 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_192 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_384 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_383 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_48 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_192 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_191 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_190 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_189 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module bit4_12 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_48 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_47 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_46 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_45 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n6), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n6), .Z(sum4[0]) );
  CND2X1 U3 ( .A(c_out400), .B(n6), .Z(n1) );
  CND2X1 U4 ( .A(c_out401), .B(c_in4), .Z(n2) );
  CND2X2 U5 ( .A(n1), .B(n2), .Z(n3) );
  CMX2X1 U6 ( .A0(s43[1]), .A1(s44[1]), .S(n3), .Z(sum4[3]) );
  CMX2X1 U7 ( .A0(s43[0]), .A1(s44[0]), .S(n3), .Z(sum4[2]) );
  CIVX1 U10 ( .A(c_out411), .Z(n4) );
  CIVX1 U11 ( .A(c_out410), .Z(n5) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(n3), .Z(c_out4) );
  CIVX2 U13 ( .A(c_in4), .Z(n6) );
endmodule


module bit8_3 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_12 A81 ( .sum4(s81), .c_out4(c_out800), .a4({a8[3:2], n2, a8[0]}), .b4(
        b8[3:0]), .c_in4(1'b0) );
  bit4_11 A82 ( .sum4(s82), .c_out4(c_out801), .a4({a8[3:2], n2, a8[0]}), .b4(
        b8[3:0]), .c_in4(1'b1) );
  bit4_10 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_9 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CND2X2 U3 ( .A(c_out810), .B(n1), .Z(n5) );
  CND2IX2 U4 ( .B(n3), .A(c_out811), .Z(n4) );
  CND2X4 U5 ( .A(n5), .B(n4), .Z(c_out8) );
  CMXI2X1 U6 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CNIVX4 U7 ( .A(a8[1]), .Z(n2) );
  CIVX1 U8 ( .A(n1), .Z(n6) );
  CMX2XL U9 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2XL U10 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2XL U11 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2XL U12 ( .A0(s81[0]), .A1(s82[0]), .S(c_in8), .Z(sum8[0]) );
  CMX2X1 U13 ( .A0(s83[3]), .A1(s84[3]), .S(n6), .Z(sum8[7]) );
  CMX2X1 U14 ( .A0(s83[2]), .A1(s84[2]), .S(n6), .Z(sum8[6]) );
  CMX2X1 U15 ( .A0(s83[0]), .A1(s84[0]), .S(n6), .Z(sum8[4]) );
  CMX2X1 U16 ( .A0(s83[1]), .A1(s84[1]), .S(n6), .Z(sum8[5]) );
  CMXI2X1 U17 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n3) );
endmodule


module Add_half_385 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_386 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_193 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_386 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_385 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_387 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_388 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_194 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_388 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_387 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_389 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(n1), .Z(sum) );
endmodule


module Add_half_390 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_195 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_390 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_389 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_391 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_392 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX1 U1 ( .A(a), .B(n1), .Z(sum) );
  CIVX20 U2 ( .A(b), .Z(n1) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_196 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_392 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_391 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_49 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_196 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_195 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_194 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_193 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CIVX1 U3 ( .A(n1), .Z(n2) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_393 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_394 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_197 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_394 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_393 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_395 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_396 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_198 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_396 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_395 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_397 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_398 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_199 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_398 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_397 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_399 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_400 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_200 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_400 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_399 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_50 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_200 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_199 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_198 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_197 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMXI2XL U3 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX1 U4 ( .A(n1), .Z(n2) );
  CIVX1 U5 ( .A(s3), .Z(n4) );
  CMX2X1 U6 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(s4), .Z(n3) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_401 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_402 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_201 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_402 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_401 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_403 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_404 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_202 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_404 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_403 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_405 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_406 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_203 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_406 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_405 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_407 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_408 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_204 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_408 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_407 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_51 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_204 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_203 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_202 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_201 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module Add_half_409 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_410 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_205 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_410 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_409 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_411 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_412 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_206 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_412 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_411 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_413 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_414 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_207 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_414 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_413 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_415 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_416 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_208 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_416 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_415 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_52 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_208 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_207 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_206 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_205 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module bit4_13 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_52 A41 ( .sum2(s41), .c_out2(c_out400), .a2({n1, a4[0]}), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_51 A42 ( .sum2(s42), .c_out2(c_out401), .a2({n1, a4[0]}), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_50 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_49 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n5), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n5), .Z(sum4[0]) );
  CNIVX2 U3 ( .A(a4[1]), .Z(n1) );
  CIVX1 U4 ( .A(c_out411), .Z(n3) );
  CMX2XL U5 ( .A0(s43[1]), .A1(s44[1]), .S(n2), .Z(sum4[3]) );
  CMX2XL U6 ( .A0(s43[0]), .A1(s44[0]), .S(n2), .Z(sum4[2]) );
  CMX2X1 U7 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CIVX2 U10 ( .A(c_out410), .Z(n4) );
  CMXI2X1 U11 ( .A0(n4), .A1(n3), .S(n2), .Z(c_out4) );
  CIVX2 U12 ( .A(c_in4), .Z(n5) );
endmodule


module Add_half_417 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_418 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_209 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_418 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_417 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_419 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_420 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_210 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_420 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_419 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_421 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_422 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_211 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_422 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_421 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_423 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_424 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_212 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_424 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_423 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_53 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_212 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_211 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_210 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_209 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CND2X1 U3 ( .A(c_out00), .B(n1), .Z(n2) );
  CND2X1 U4 ( .A(c_out01), .B(c_in2), .Z(n3) );
  CND2X2 U5 ( .A(n2), .B(n3), .Z(n4) );
  CIVX2 U6 ( .A(c_in2), .Z(n1) );
  CMXI2XL U8 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CMX2X1 U9 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_425 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_426 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_213 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_426 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_425 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_427 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_428 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_214 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_428 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_427 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_429 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(n2) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U4 ( .A(b), .B(n2), .Z(sum) );
endmodule


module Add_half_430 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_215 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_430 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_429 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_431 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_432 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_216 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_432 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_431 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_54 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_216 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_215 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_214 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_213 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n1), .Z(sum2[0]) );
  CND2X1 U3 ( .A(c_out00), .B(n1), .Z(n2) );
  CND2X2 U4 ( .A(c_out01), .B(c_in2), .Z(n3) );
  CND2X2 U5 ( .A(n2), .B(n3), .Z(n4) );
  CIVX2 U6 ( .A(c_in2), .Z(n1) );
  CMXI2XL U8 ( .A0(n8), .A1(n7), .S(n4), .Z(sum2[1]) );
  CIVX1 U9 ( .A(s3), .Z(n8) );
  CIVX2 U10 ( .A(c_out10), .Z(n6) );
  CIVX2 U11 ( .A(c_out11), .Z(n5) );
  CMXI2X1 U12 ( .A0(n6), .A1(n5), .S(n4), .Z(c_out2) );
  CIVX2 U13 ( .A(s4), .Z(n7) );
endmodule


module Add_half_433 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_434 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_217 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_434 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_433 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_435 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_436 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_218 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_436 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_435 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_437 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_438 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_219 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_438 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_437 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_439 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_440 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_220 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_440 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_439 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_55 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_220 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_219 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_218 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_217 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(n1), .Z(n4) );
  CMXI2XL U4 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_441 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_442 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_221 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_442 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_441 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_443 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_444 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_222 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_444 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_443 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_445 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_446 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_223 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_446 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_445 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_447 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_448 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_224 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_448 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_447 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_56 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_224 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_223 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_222 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_221 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2XL U4 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CIVX1 U5 ( .A(c_out11), .Z(n2) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module bit4_14 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_56 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_55 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_54 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_53 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMX2XL U4 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2XL U5 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2X1 U6 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_449 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_450 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_225 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_450 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_449 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_451 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_452 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_226 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_452 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_451 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_453 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_454 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_227 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_454 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_453 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_455 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_456 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_228 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_456 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_455 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_57 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_228 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_227 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_226 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_225 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_457 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_458 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_229 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_458 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_457 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_459 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_460 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_230 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_460 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_459 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_461 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_462 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_231 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_462 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_461 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_463 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_464 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_232 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_464 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_463 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_58 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_232 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_231 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_230 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_229 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_465 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_466 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_233 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_466 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_465 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_467 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_468 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_234 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_468 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_467 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_469 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_470 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_235 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_470 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_469 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_471 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_472 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_236 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_472 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_471 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_59 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_236 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_235 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_234 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_233 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n5) );
  CIVX2 U5 ( .A(c_out10), .Z(n2) );
  CIVX2 U8 ( .A(c_out11), .Z(n1) );
  CMXI2X1 U9 ( .A0(n2), .A1(n1), .S(n5), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n4) );
endmodule


module Add_half_473 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_474 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_237 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_474 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_473 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_475 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_476 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_238 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_476 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_475 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_477 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_478 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_239 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_478 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_477 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_479 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_480 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_240 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_480 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_479 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_60 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_240 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_239 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_238 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_237 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n5) );
  CIVX2 U5 ( .A(c_out10), .Z(n2) );
  CIVX2 U8 ( .A(c_out11), .Z(n1) );
  CMXI2X1 U9 ( .A0(n2), .A1(n1), .S(n5), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n4) );
endmodule


module bit4_15 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_60 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_59 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_58 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_57 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n8), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n8), .Z(sum4[0]) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum4[2]) );
  CMXI2XL U4 ( .A0(n7), .A1(n6), .S(n1), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX1 U6 ( .A(c_out411), .Z(n2) );
  CIVX1 U7 ( .A(c_out410), .Z(n3) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out4) );
  CIVX2 U11 ( .A(s43[0]), .Z(n5) );
  CIVX2 U12 ( .A(s44[0]), .Z(n4) );
  CIVX2 U13 ( .A(s43[1]), .Z(n7) );
  CIVX2 U14 ( .A(s44[1]), .Z(n6) );
  CIVX2 U15 ( .A(c_in4), .Z(n8) );
endmodule


module Add_half_481 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_482 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_241 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_482 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_481 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_483 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_484 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_242 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_484 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_483 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_485 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_486 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_243 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_486 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_485 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_487 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_488 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_244 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_488 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_487 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_61 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_244 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_243 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_242 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_241 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_489 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_490 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_245 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_490 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_489 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_491 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_492 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_246 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_492 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_491 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_493 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_494 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_247 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_494 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_493 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_495 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_496 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_248 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_496 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_495 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_62 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_248 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_247 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_246 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_245 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_497 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_498 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_249 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_498 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_497 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_499 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_500 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_250 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_500 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_499 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_501 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_502 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_251 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_502 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_501 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_503 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_504 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_252 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_504 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_503 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_63 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_252 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_251 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_250 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_249 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n5) );
  CIVX2 U5 ( .A(c_out10), .Z(n2) );
  CIVX2 U8 ( .A(c_out11), .Z(n1) );
  CMXI2X1 U9 ( .A0(n2), .A1(n1), .S(n5), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n4) );
endmodule


module Add_half_505 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_506 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_253 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_506 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_505 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_507 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_508 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_254 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_508 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_507 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_509 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_510 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_255 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_510 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_509 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_511 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_512 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_256 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_512 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_511 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_64 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_256 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_255 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_254 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_253 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n5) );
  CIVX2 U5 ( .A(c_out10), .Z(n2) );
  CIVX2 U8 ( .A(c_out11), .Z(n1) );
  CMXI2X1 U9 ( .A0(n2), .A1(n1), .S(n5), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n4) );
endmodule


module bit4_16 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_64 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_63 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_62 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_61 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n8), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n8), .Z(sum4[0]) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum4[2]) );
  CMXI2XL U4 ( .A0(n7), .A1(n6), .S(n1), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX1 U6 ( .A(c_out411), .Z(n2) );
  CIVX1 U7 ( .A(c_out410), .Z(n3) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out4) );
  CIVX2 U11 ( .A(s43[0]), .Z(n5) );
  CIVX2 U12 ( .A(s44[0]), .Z(n4) );
  CIVX2 U13 ( .A(s43[1]), .Z(n7) );
  CIVX2 U14 ( .A(s44[1]), .Z(n6) );
  CIVX2 U15 ( .A(c_in4), .Z(n8) );
endmodule


module bit8_4 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_16 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_15 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_14 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_13 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n3), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n3), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n3), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n3), .Z(sum8[0]) );
  CMXI2X1 U3 ( .A0(c_out810), .A1(c_out811), .S(n2), .Z(n1) );
  CIVX2 U4 ( .A(n1), .Z(c_out8) );
  CMX2XL U5 ( .A0(s83[2]), .A1(s84[2]), .S(n2), .Z(sum8[6]) );
  CMX2XL U6 ( .A0(s83[3]), .A1(s84[3]), .S(n2), .Z(sum8[7]) );
  CMX2XL U7 ( .A0(s83[1]), .A1(s84[1]), .S(n2), .Z(sum8[5]) );
  CMX2XL U8 ( .A0(s83[0]), .A1(s84[0]), .S(n2), .Z(sum8[4]) );
  CMX2X1 U9 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n2) );
  CIVX2 U14 ( .A(c_in8), .Z(n3) );
endmodule


module bit32_1 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   c1, c2, c3, n1, n2, n3, n4, n5, n6, n7;

  bit8_4 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8(a32[7:0]), .b8(b32[7:0]), 
        .c_in8(c_in32) );
  bit8_3 A322 ( .sum8(sum32[15:8]), .c_out8(c2), .a8({a32[15], n5, a32[13:8]}), 
        .b8({b32[15:14], n1, b32[12:8]}), .c_in8(c1) );
  bit8_2 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8({a32[23], n3, a32[21:16]}), .b8(b32[23:16]), .c_in8(c2) );
  bit8_1 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8({a32[31:26], n7, 
        a32[24]}), .b8(b32[31:24]), .c_in8(c3) );
  CNIVX3 U1 ( .A(b32[13]), .Z(n1) );
  CIVX4 U2 ( .A(a32[25]), .Z(n6) );
  CIVX8 U3 ( .A(n6), .Z(n7) );
  CIVX1 U4 ( .A(a32[22]), .Z(n2) );
  CIVX4 U5 ( .A(n2), .Z(n3) );
  CIVX1 U6 ( .A(a32[14]), .Z(n4) );
  CIVX4 U7 ( .A(n4), .Z(n5) );
endmodule


module Add_half_513 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_514 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_257 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_514 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_513 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_515 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_516 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_258 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_516 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_515 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_517 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_518 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_259 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_518 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_517 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_519 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_520 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_260 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_520 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_519 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_65 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_260 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_259 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_258 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_257 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(s3), .Z(n3) );
  CIVX2 U7 ( .A(s4), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(sum2[1]) );
endmodule


module Add_half_521 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n1) );
  CENX1 U3 ( .A(a), .B(n1), .Z(sum) );
endmodule


module Add_half_522 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_261 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_522 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_521 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_523 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_524 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_262 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_524 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_523 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_525 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_526 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_263 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_526 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_525 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_527 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_528 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_264 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_528 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_527 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_66 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_264 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_263 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_262 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_261 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_529 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_530 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_265 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_530 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_529 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_531 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_532 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_266 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_532 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_531 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_533 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_534 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_267 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_534 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_533 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_535 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_536 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_268 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_536 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_535 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_67 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_268 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_267 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_266 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_265 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s2), .Z(n4) );
  CIVX1 U4 ( .A(s1), .Z(n5) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n6) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_537 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_538 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_269 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_538 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_537 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_539 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_540 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_270 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_540 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_539 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_541 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_542 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_271 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_542 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_541 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_543 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_544 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_272 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_544 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_543 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_68 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_272 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_271 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_270 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_269 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_17 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_68 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_67 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_66 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_65 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMX2X1 U4 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U7 ( .A(s41[1]), .Z(n3) );
  CIVX2 U8 ( .A(s42[1]), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U10 ( .A(s43[0]), .Z(n5) );
  CIVX2 U11 ( .A(s44[0]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(n1), .Z(sum4[2]) );
endmodule


module Add_half_545 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_546 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_273 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_546 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_545 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_547 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_548 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_274 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_548 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_547 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_549 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_550 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_275 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_550 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_549 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_551 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_552 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_276 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_552 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_551 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_69 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_276 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_275 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_274 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_273 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CIVX2 U7 ( .A(s1), .Z(n3) );
  CIVX2 U8 ( .A(s2), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_553 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_554 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_277 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_554 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_553 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_555 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_556 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_278 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_556 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_555 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_557 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_558 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_279 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_558 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_557 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_559 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_560 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_280 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_560 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_559 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_70 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_280 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_279 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_278 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_277 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_561 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_562 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_281 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_562 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_561 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_563 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_564 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_282 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_564 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_563 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_565 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_566 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_283 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_566 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_565 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_567 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_568 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_284 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_568 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_567 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_71 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_284 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_283 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_282 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_281 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2XL U4 ( .A0(n7), .A1(n6), .S(n5), .Z(sum2[1]) );
  CIVX1 U5 ( .A(n2), .Z(n5) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out10), .Z(n4) );
  CIVX2 U9 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(n5), .Z(c_out2) );
  CIVX2 U11 ( .A(s3), .Z(n7) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
endmodule


module Add_half_569 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_570 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_285 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_570 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_569 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_571 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_572 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_286 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_572 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_571 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_573 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_574 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_287 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_574 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_573 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_575 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_576 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_288 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_576 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_575 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_72 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_288 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_287 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_286 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_285 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(n1), .Z(n4) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_18 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_72 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_71 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_70 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_69 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n1), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CMX2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMX2X1 U6 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2X1 U7 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U8 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX1 U9 ( .A(s43[1]), .Z(n3) );
  CIVX2 U10 ( .A(s44[1]), .Z(n2) );
endmodule


module Add_half_577 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_578 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_289 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_578 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_577 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_579 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_580 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_290 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_580 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_579 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_581 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_582 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_291 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_582 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_581 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_583 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_584 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2XL U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX2 U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_292 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_584 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_583 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_73 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8, n9;

  Add_full_292 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_291 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_290 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_289 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2X2 U3 ( .A(c_out10), .B(n1), .Z(n2) );
  CND2X2 U4 ( .A(c_out11), .B(n7), .Z(n3) );
  CND2X2 U5 ( .A(n2), .B(n3), .Z(c_out2) );
  CIVX2 U6 ( .A(n7), .Z(n1) );
  CMXI2XL U7 ( .A0(n9), .A1(n8), .S(n7), .Z(sum2[1]) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n4) );
  CIVX2 U9 ( .A(n4), .Z(n7) );
  CIVX2 U10 ( .A(s1), .Z(n6) );
  CIVX2 U11 ( .A(s2), .Z(n5) );
  CMXI2X1 U12 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U13 ( .A(s3), .Z(n9) );
  CIVX2 U14 ( .A(s4), .Z(n8) );
endmodule


module Add_half_585 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_586 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_293 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_586 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_585 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_587 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_588 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_294 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_588 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_587 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_589 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_590 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_295 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_590 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_589 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_591 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_592 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_296 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_592 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_591 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_74 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_296 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_295 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_294 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_293 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n4), .S(n2), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_in2), .Z(n1) );
  CMX2X1 U5 ( .A0(c_out11), .A1(c_out10), .S(n2), .Z(c_out2) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(s3), .Z(n4) );
  CIVX2 U9 ( .A(s4), .Z(n3) );
endmodule


module Add_half_593 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_594 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_297 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_594 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_593 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_595 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_596 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_298 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_596 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_595 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_597 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_598 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_299 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_598 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_597 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_599 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_600 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_300 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_600 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_599 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_75 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_300 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_299 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_298 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_297 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s2), .Z(n5) );
  CIVX1 U4 ( .A(s1), .Z(n6) );
  CMX2XL U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U6 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CIVX2 U7 ( .A(c_out10), .Z(n4) );
  CIVX2 U8 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMXI2X1 U10 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n1), .Z(sum2[1]) );
endmodule


module Add_half_601 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_602 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_301 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_602 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_601 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_603 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_604 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_302 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_604 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_603 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_605 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_606 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_303 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_606 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_605 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX1 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_607 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_608 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_304 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_608 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_607 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_76 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_304 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_303 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_302 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_301 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMX2XL U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U5 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out10), .Z(n4) );
  CIVX2 U9 ( .A(c_out11), .Z(n3) );
endmodule


module bit4_19 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_76 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_75 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_74 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_73 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(n3), .Z(n1) );
  CIVX2 U4 ( .A(c_in4), .Z(n2) );
  CIVX1 U5 ( .A(s44[1]), .Z(n6) );
  CIVX1 U6 ( .A(s43[1]), .Z(n7) );
  CMXI2X1 U7 ( .A0(c_out401), .A1(c_out400), .S(n2), .Z(n3) );
  CMXI2XL U8 ( .A0(n7), .A1(n6), .S(n1), .Z(sum4[3]) );
  CMX2XL U9 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2X1 U10 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U11 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U12 ( .A(c_out410), .Z(n5) );
  CIVX2 U13 ( .A(c_out411), .Z(n4) );
  CMXI2X1 U14 ( .A0(n5), .A1(n4), .S(n1), .Z(c_out4) );
endmodule


module Add_half_609 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_610 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_305 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_610 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_609 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_611 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_612 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_306 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_612 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_611 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_613 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_614 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_307 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_614 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_613 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_615 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_616 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_308 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_616 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_615 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_77 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1;

  Add_full_308 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_307 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_306 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_305 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_617 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_618 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_309 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_618 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_617 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_619 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_620 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_310 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_620 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_619 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_621 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_622 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_311 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_622 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_621 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_623 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_624 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_312 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_624 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_623 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_78 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_312 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_311 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_310 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_309 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2X2 U3 ( .A(c_out10), .B(n1), .Z(n2) );
  CND2X2 U4 ( .A(c_out11), .B(n5), .Z(n3) );
  CND2X2 U5 ( .A(n2), .B(n3), .Z(c_out2) );
  CIVX2 U6 ( .A(n5), .Z(n1) );
  CMXI2XL U7 ( .A0(n7), .A1(n6), .S(n5), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n4) );
  CIVX2 U10 ( .A(n4), .Z(n5) );
  CIVX2 U11 ( .A(s3), .Z(n7) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
endmodule


module Add_half_625 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_626 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_313 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_626 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_625 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_627 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_628 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_314 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_628 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_627 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_629 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_630 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_315 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_630 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_629 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_631 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_632 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_316 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_632 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_631 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_79 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_316 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_315 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_314 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_313 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(n1), .Z(n4) );
  CMXI2X1 U4 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out10), .Z(n3) );
  CIVX2 U9 ( .A(c_out11), .Z(n2) );
endmodule


module Add_half_633 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_634 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_317 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_634 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_633 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_635 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_636 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_318 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_636 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_635 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_637 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_638 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_319 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_638 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_637 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_639 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_640 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_320 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_640 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_639 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_80 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_320 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_319 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_318 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_317 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(n1), .Z(n4) );
  CMXI2X1 U4 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out10), .Z(n3) );
  CIVX2 U9 ( .A(c_out11), .Z(n2) );
endmodule


module bit4_20 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_80 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_79 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_78 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_77 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(c_in4), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out401), .A1(c_out400), .S(n1), .Z(n2) );
  CIVX2 U5 ( .A(c_out410), .Z(n4) );
  CIVX1 U6 ( .A(s43[0]), .Z(n6) );
  CMXI2XL U7 ( .A0(n6), .A1(n5), .S(n7), .Z(sum4[2]) );
  CMX2XL U8 ( .A0(s43[1]), .A1(s44[1]), .S(n7), .Z(sum4[3]) );
  CMX2X1 U9 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U10 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U11 ( .A(c_out411), .Z(n3) );
  CIVX2 U12 ( .A(n2), .Z(n7) );
  CMXI2X1 U13 ( .A0(n4), .A1(n3), .S(n7), .Z(c_out4) );
  CIVX2 U14 ( .A(s44[0]), .Z(n5) );
endmodule


module bit8_5 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   n19, n20, c_out800, c_out801, c_out810, c_out811, n2, n3, n4, n5, n6,
         n7, n8, n9, n11, n12, n13, n14, n15, n16, n17, n18;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_20 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4({b8[3:2], n12, 
        b8[0]}), .c_in4(1'b0) );
  bit4_19 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4({b8[3:2], n12, 
        b8[0]}), .c_in4(1'b1) );
  bit4_18 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_17 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CNIVX4 U3 ( .A(n19), .Z(sum8[1]) );
  CMX2X2 U4 ( .A0(s83[3]), .A1(s84[3]), .S(n3), .Z(sum8[7]) );
  CIVX2 U5 ( .A(n20), .Z(n9) );
  CMXI2X1 U6 ( .A0(n15), .A1(n16), .S(n6), .Z(n20) );
  CIVX2 U7 ( .A(c_in8), .Z(n6) );
  CIVXL U8 ( .A(n8), .Z(n2) );
  CIVX1 U9 ( .A(n2), .Z(n3) );
  CMX2XL U10 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(n19) );
  CND2X1 U11 ( .A(s83[2]), .B(n2), .Z(n4) );
  CND2XL U12 ( .A(s84[2]), .B(n8), .Z(n5) );
  CND2X2 U13 ( .A(n4), .B(n5), .Z(sum8[6]) );
  CIVX8 U14 ( .A(n9), .Z(sum8[0]) );
  CIVX1 U15 ( .A(n6), .Z(n7) );
  CIVX1 U16 ( .A(b8[1]), .Z(n11) );
  CMX2X2 U17 ( .A0(s81[3]), .A1(s82[3]), .S(n7), .Z(sum8[3]) );
  CMX2X2 U18 ( .A0(s81[2]), .A1(s82[2]), .S(n7), .Z(sum8[2]) );
  CMX2X2 U19 ( .A0(s83[1]), .A1(s84[1]), .S(n8), .Z(sum8[5]) );
  CMX2X2 U20 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n8) );
  CIVX1 U21 ( .A(s84[0]), .Z(n17) );
  CIVX4 U22 ( .A(n11), .Z(n12) );
  CMXI2XL U23 ( .A0(n14), .A1(n13), .S(n3), .Z(c_out8) );
  CMXI2X1 U24 ( .A0(n18), .A1(n17), .S(n8), .Z(sum8[4]) );
  CIVX2 U25 ( .A(c_out810), .Z(n14) );
  CIVX2 U26 ( .A(c_out811), .Z(n13) );
  CIVX2 U27 ( .A(s81[0]), .Z(n16) );
  CIVX2 U28 ( .A(s82[0]), .Z(n15) );
  CIVX2 U29 ( .A(s83[0]), .Z(n18) );
endmodule


module Add_half_641 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_642 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_321 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_642 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_641 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_643 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_644 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_322 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_644 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_643 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_645 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_646 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_323 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_646 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_645 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_647 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_648 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_324 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_648 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_647 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_81 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_324 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_323 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_322 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_321 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_649 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_650 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_325 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_650 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_649 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_651 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_652 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_326 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_652 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_651 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_653 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_654 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_327 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_654 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_653 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_655 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_656 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_328 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_656 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_655 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_82 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_328 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_327 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_326 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_325 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_657 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_658 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_329 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_658 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_657 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_659 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_660 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_330 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_660 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_659 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_661 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_662 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_331 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_662 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_661 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_663 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_664 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_332 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_664 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_663 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_83 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_332 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_331 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_330 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_329 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_665 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_666 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_333 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_666 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_665 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_667 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_668 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_334 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_668 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_667 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_669 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_670 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_335 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_670 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_669 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_671 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_672 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_336 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_672 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_671 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_84 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_336 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_335 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_334 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_333 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s2), .Z(n4) );
  CIVX1 U4 ( .A(s1), .Z(n5) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n6) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module bit4_21 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_84 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_83 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_82 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_81 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
  CIVXL U4 ( .A(c_out411), .Z(n2) );
  CIVX2 U5 ( .A(c_out410), .Z(n3) );
  CMX2XL U6 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2XL U7 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U8 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U9 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMXI2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U11 ( .A(n1), .Z(n4) );
endmodule


module Add_half_673 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_674 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_337 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_674 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_673 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_675 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_676 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_338 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_676 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_675 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_677 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_678 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_339 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_678 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_677 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_679 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_680 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_340 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_680 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_679 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_85 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_340 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_339 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_338 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_337 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_681 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_682 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_341 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_682 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_681 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_683 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_684 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_342 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_684 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_683 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_685 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_686 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_343 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_686 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_685 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_687 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_688 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_344 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_688 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_687 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_86 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1;

  Add_full_344 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_343 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_342 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_341 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_689 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_690 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_345 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_690 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_689 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_691 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_692 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_346 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_692 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_691 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_693 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_694 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_347 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_694 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_693 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_695 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_696 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVX1 U1 ( .A(b), .Z(n2) );
  CND2X1 U2 ( .A(a), .B(n2), .Z(n3) );
  CIVX1 U3 ( .A(a), .Z(n1) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CND2X1 U5 ( .A(n1), .B(b), .Z(n4) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_348 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_696 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_695 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_87 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_348 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_347 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_346 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_345 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U4 ( .A(n1), .Z(n4) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_697 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_698 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_349 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_698 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_697 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_699 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_700 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_350 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_700 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_699 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_701 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_702 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_351 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_702 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_701 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_703 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_704 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(n2), .B(a), .Z(n3) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CIVX1 U3 ( .A(a), .Z(n1) );
  CND2X1 U4 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U5 ( .A(n3), .B(n4), .Z(sum) );
  CAN2XL U6 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_352 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_704 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_703 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_88 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_352 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_351 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_350 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_349 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n2) );
  CIVX1 U5 ( .A(c_out11), .Z(n4) );
  CMX2X1 U6 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVXL U7 ( .A(n2), .Z(n1) );
  CIVXL U8 ( .A(n1), .Z(n6) );
  CMX2X1 U9 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U10 ( .A(c_out10), .Z(n5) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(n2), .Z(c_out2) );
endmodule


module bit4_22 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_88 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_87 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_86 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_85 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n10), .A1(n11), .S(n1), .Z(sum4[3]) );
  CIVXL U4 ( .A(n9), .Z(n1) );
  CIVX1 U5 ( .A(s41[1]), .Z(n6) );
  CIVX1 U6 ( .A(s42[0]), .Z(n3) );
  CMXI2XL U7 ( .A0(n8), .A1(n7), .S(n9), .Z(sum4[2]) );
  CMX2X1 U8 ( .A0(c_out410), .A1(c_out411), .S(n9), .Z(c_out4) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CIVX2 U10 ( .A(n2), .Z(n9) );
  CIVX2 U11 ( .A(s41[0]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n4), .A1(n3), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U13 ( .A(s42[1]), .Z(n5) );
  CMXI2X1 U14 ( .A0(n6), .A1(n5), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U15 ( .A(s43[0]), .Z(n8) );
  CIVX2 U16 ( .A(s44[0]), .Z(n7) );
  CIVX2 U17 ( .A(s43[1]), .Z(n11) );
  CIVX2 U18 ( .A(s44[1]), .Z(n10) );
endmodule


module Add_half_705 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_706 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_353 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_706 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_705 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_707 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_708 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_354 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_708 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_707 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_709 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_710 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_355 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_710 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_709 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_711 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_712 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_356 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_712 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_711 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_89 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_356 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_355 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_354 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_353 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n7), .A1(n6), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n7) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
endmodule


module Add_half_713 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_714 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_357 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_714 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_713 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_715 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_716 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_358 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_716 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_715 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_717 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_718 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_359 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_718 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_717 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_719 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_720 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_360 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_720 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_719 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_90 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_360 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_359 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_358 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_357 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
endmodule


module Add_half_721 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_722 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_361 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_722 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_721 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_723 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_724 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_362 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_724 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_723 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_725 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_726 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_363 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_726 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_725 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_727 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_728 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_364 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_728 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_727 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_91 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_364 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_363 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_362 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_361 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_729 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_730 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_365 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_730 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_729 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_731 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_732 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_366 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_732 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_731 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_733 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_734 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_367 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_734 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_733 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_735 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_736 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_368 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_736 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_735 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_92 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_368 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_367 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_366 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_365 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_23 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_92 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_91 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_90 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_89 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n6), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n6), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n6) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out4) );
  CIVX2 U11 ( .A(s41[1]), .Z(n5) );
  CIVX2 U12 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
endmodule


module Add_half_737 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_738 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_369 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_738 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_737 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_739 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_740 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_370 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_740 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_739 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_741 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_742 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_371 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_742 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_741 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_743 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_744 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_372 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_744 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_743 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_93 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_372 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_371 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_370 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_369 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_745 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_746 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_373 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_746 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_745 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_747 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_748 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_374 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_748 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_747 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_749 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_750 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_375 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_750 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_749 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_751 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_752 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_376 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_752 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_751 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_94 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_376 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_375 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_374 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_373 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_753 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_754 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_377 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_754 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_753 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_755 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_756 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_378 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_756 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_755 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_757 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_758 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_379 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_758 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_757 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_759 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_760 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_380 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_760 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_759 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_95 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_380 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_379 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_378 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_377 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_761 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_762 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_381 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_762 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_761 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_763 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_764 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_382 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_764 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_763 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_765 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_766 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_383 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_766 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_765 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_767 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_768 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_384 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_768 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_767 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_96 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_384 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_383 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_382 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_381 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_24 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_96 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_95 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_94 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_93 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX1 U4 ( .A(c_out411), .Z(n2) );
  CIVX2 U5 ( .A(n1), .Z(n8) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CMXI2X1 U7 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U9 ( .A(s41[0]), .Z(n5) );
  CIVX2 U10 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U12 ( .A(s43[0]), .Z(n7) );
  CIVX2 U13 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX2 U15 ( .A(s43[1]), .Z(n10) );
  CIVX2 U16 ( .A(s44[1]), .Z(n9) );
  CMXI2X1 U17 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
endmodule


module bit8_6 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   n14, c_out800, c_out801, c_out810, c_out811, n1, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_24 A81 ( .sum4(s81), .c_out4(c_out800), .a4({a8[3:1], n3}), .b4(b8[3:0]), .c_in4(1'b0) );
  bit4_23 A82 ( .sum4(s82), .c_out4(c_out801), .a4({a8[3:1], n3}), .b4(b8[3:0]), .c_in4(1'b1) );
  bit4_22 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_21 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X2 U3 ( .A0(s83[2]), .A1(s84[2]), .S(n13), .Z(sum8[6]) );
  CIVX2 U4 ( .A(n14), .Z(n1) );
  CIVX4 U5 ( .A(n1), .Z(sum8[1]) );
  CMXI2X1 U6 ( .A0(n8), .A1(n7), .S(n5), .Z(n14) );
  CIVX1 U7 ( .A(n6), .Z(n13) );
  CMXI2X1 U8 ( .A0(n10), .A1(n9), .S(n13), .Z(sum8[4]) );
  CMX2X2 U9 ( .A0(s81[0]), .A1(s82[0]), .S(c_in8), .Z(sum8[0]) );
  CNIVX4 U10 ( .A(a8[0]), .Z(n3) );
  CMX2X1 U11 ( .A0(c_out811), .A1(c_out810), .S(n6), .Z(c_out8) );
  CIVX1 U12 ( .A(s83[1]), .Z(n12) );
  CMX2X2 U13 ( .A0(s81[2]), .A1(s82[2]), .S(n5), .Z(sum8[2]) );
  CIVX2 U14 ( .A(n4), .Z(n5) );
  CIVXL U15 ( .A(c_in8), .Z(n4) );
  CMX2XL U16 ( .A0(s83[3]), .A1(s84[3]), .S(n13), .Z(sum8[7]) );
  CMX2X1 U17 ( .A0(s81[3]), .A1(s82[3]), .S(n5), .Z(sum8[3]) );
  CMXI2X2 U18 ( .A0(n12), .A1(n11), .S(n13), .Z(sum8[5]) );
  CMXI2X1 U19 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n6) );
  CIVX2 U20 ( .A(s81[1]), .Z(n8) );
  CIVX2 U21 ( .A(s82[1]), .Z(n7) );
  CIVX2 U22 ( .A(s83[0]), .Z(n10) );
  CIVX2 U23 ( .A(s84[0]), .Z(n9) );
  CIVX2 U24 ( .A(s84[1]), .Z(n11) );
endmodule


module Add_half_769 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_770 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_385 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_770 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_769 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_771 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_772 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_386 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_772 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_771 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_773 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_774 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_387 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_774 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_773 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_775 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_776 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_388 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_776 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_775 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_97 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_388 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_387 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_386 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_385 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_777 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_778 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_389 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_778 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_777 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_779 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_780 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_390 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_780 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_779 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_781 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_782 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_391 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_782 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_781 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_783 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_784 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_392 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_784 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_783 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_98 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_392 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_391 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_390 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_389 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_785 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_786 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_393 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_786 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_785 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_787 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_788 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_394 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_788 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_787 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_789 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_790 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_395 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_790 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_789 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_791 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_792 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_396 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_792 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_791 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_99 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_396 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_395 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_394 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_393 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_793 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_794 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_397 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_794 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_793 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_795 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_796 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_398 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_796 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_795 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_797 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_798 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_399 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_798 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_797 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_799 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_800 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_400 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_800 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_799 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_100 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_400 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_399 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_398 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_397 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CMXI2XL U4 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n4) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module bit4_25 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_100 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_99 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_98 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_97 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U4 ( .A0(c_out410), .A1(c_out411), .S(n4), .Z(c_out4) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CIVX2 U8 ( .A(s41[0]), .Z(n3) );
  CIVX2 U9 ( .A(s42[0]), .Z(n2) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U11 ( .A(s43[1]), .Z(n6) );
  CIVX2 U12 ( .A(s44[1]), .Z(n5) );
  CMXI2X1 U13 ( .A0(n6), .A1(n5), .S(n4), .Z(sum4[3]) );
endmodule


module Add_half_801 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_802 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_401 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_802 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_801 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_803 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_804 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_402 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_804 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_803 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_805 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_806 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_403 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_806 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_805 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_807 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_808 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVXL U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_404 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_808 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_807 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_101 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_404 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_403 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_402 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_401 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U7 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_809 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_810 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_405 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_810 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_809 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_811 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_812 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_406 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_812 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_811 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_813 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_814 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_407 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_814 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_813 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_815 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_816 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_408 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_816 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_815 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_102 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_408 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_407 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_406 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_405 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_817 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_818 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_409 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_818 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_817 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_819 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_820 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_410 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_820 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_819 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_821 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_822 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_411 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_822 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_821 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_823 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_824 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_412 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_824 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_823 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_103 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_412 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_411 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_410 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_409 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_825 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_826 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_413 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_826 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_825 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_827 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_828 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_414 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_828 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_827 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_829 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_830 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_415 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_830 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_829 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_831 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_832 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_416 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_832 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_831 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_104 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_416 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_415 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_414 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_413 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_26 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_104 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_103 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_102 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_101 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(s44[0]), .Z(n4) );
  CMX2XL U4 ( .A0(s43[1]), .A1(s44[1]), .S(n6), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n6) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out4) );
  CIVX2 U12 ( .A(s43[0]), .Z(n5) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(n6), .Z(sum4[2]) );
endmodule


module Add_half_833 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_834 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_417 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_834 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_833 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_835 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_836 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_418 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_836 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_835 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_837 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_838 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_419 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_838 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_837 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_839 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_840 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_420 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_840 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_839 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_105 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_420 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_419 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_418 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_417 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(s2), .Z(n2) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CIVX2 U7 ( .A(s1), .Z(n3) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_841 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_842 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_421 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_842 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_841 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_843 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_844 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_422 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_844 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_843 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_845 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_846 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_423 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_846 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_845 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_847 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_848 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_424 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_848 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_847 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_106 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_424 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_423 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_422 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_421 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CIVX1 U3 ( .A(s3), .Z(n4) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_849 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_850 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_425 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_850 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_849 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_851 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_852 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_426 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_852 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_851 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_853 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_854 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_427 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_854 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_853 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_855 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_856 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_428 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_856 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_855 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_107 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_428 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_427 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_426 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_425 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n3), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CIVX2 U4 ( .A(n3), .Z(n5) );
  CIVX2 U5 ( .A(c_out10), .Z(n2) );
  CIVX2 U8 ( .A(c_out11), .Z(n1) );
  CMXI2X1 U9 ( .A0(n2), .A1(n1), .S(n5), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n4) );
endmodule


module Add_half_857 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_858 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_429 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_858 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_857 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_859 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_860 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_430 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_860 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_859 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_861 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_862 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_431 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_862 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_861 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_863 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_864 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_432 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_864 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_863 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_108 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_432 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_431 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_430 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_429 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CIVX1 U4 ( .A(s3), .Z(n5) );
  CMX2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module bit4_27 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_108 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_107 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_106 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_105 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out4) );
  CIVX2 U11 ( .A(c_in4), .Z(n4) );
endmodule


module Add_half_865 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_866 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_433 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_866 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_865 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_867 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_868 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_434 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_868 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_867 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_869 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_870 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_435 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_870 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_869 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_871 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_872 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_436 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_872 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_871 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_109 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_436 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_435 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_434 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_433 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_873 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_874 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_437 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_874 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_873 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_875 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_876 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_438 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_876 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_875 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_877 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_878 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_439 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_878 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_877 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_879 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_880 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_440 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_880 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_879 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_110 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_440 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_439 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_438 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_437 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_881 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_882 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_441 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_882 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_881 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_883 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_884 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_442 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_884 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_883 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_885 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_886 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_443 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_886 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_885 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_887 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_888 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_444 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_888 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_887 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_111 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_444 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_443 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_442 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_441 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module Add_half_889 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_890 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_445 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_890 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_889 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_891 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_892 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_446 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_892 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_891 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_893 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_894 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_447 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_894 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_893 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_895 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_896 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_448 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_896 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_895 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_112 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_448 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_447 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_446 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_445 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U5 ( .A(s3), .Z(n5) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module bit4_28 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_112 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_111 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_110 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_109 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n9), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n9), .Z(sum4[0]) );
  CMXI2XL U3 ( .A0(n8), .A1(n7), .S(n6), .Z(sum4[3]) );
  CIVX1 U4 ( .A(c_out410), .Z(n3) );
  CIVX2 U5 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out4) );
  CIVX2 U11 ( .A(s43[0]), .Z(n5) );
  CIVX2 U12 ( .A(s44[0]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(n6), .Z(sum4[2]) );
  CIVX2 U14 ( .A(s43[1]), .Z(n8) );
  CIVX2 U15 ( .A(s44[1]), .Z(n7) );
  CIVX2 U16 ( .A(c_in4), .Z(n9) );
endmodule


module bit8_7 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_28 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_27 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_26 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_25 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n5), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n5), .Z(sum8[0]) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n4), .Z(sum8[5]) );
  CMX2X2 U4 ( .A0(s83[0]), .A1(s84[0]), .S(n4), .Z(sum8[4]) );
  CMX2X2 U5 ( .A0(s83[2]), .A1(s84[2]), .S(n4), .Z(sum8[6]) );
  CMX2X1 U6 ( .A0(s83[3]), .A1(s84[3]), .S(n4), .Z(sum8[7]) );
  CIVX1 U7 ( .A(s84[1]), .Z(n2) );
  CMX2X2 U8 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2X1 U9 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2X1 U10 ( .A0(c_out810), .A1(c_out811), .S(n4), .Z(c_out8) );
  CIVX2 U11 ( .A(n1), .Z(n4) );
  CMXI2X1 U14 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CIVX2 U15 ( .A(s83[1]), .Z(n3) );
  CIVX2 U16 ( .A(c_in8), .Z(n5) );
endmodule


module Add_half_897 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_898 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_449 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_898 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_897 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_899 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_900 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_450 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_900 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_899 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_901 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_902 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_451 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_902 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_901 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_903 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_904 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_452 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_904 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_903 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_113 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_452 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_451 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_450 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_449 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_905 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_906 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_453 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_906 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_905 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_907 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_908 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_454 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_908 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_907 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_909 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_910 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_455 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_910 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_909 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_911 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_912 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_456 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_912 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_911 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_114 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_456 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_455 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_454 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_453 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_913 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_914 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_457 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_914 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_913 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_915 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_916 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_458 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_916 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_915 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_917 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_918 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_459 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_918 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_917 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_919 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_920 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_460 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_920 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_919 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_115 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_460 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_459 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_458 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_457 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_921 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_922 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_461 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_922 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_921 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_923 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_924 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_462 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_924 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_923 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_925 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_926 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_463 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_926 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_925 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_927 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_928 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_464 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_928 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_927 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_116 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_464 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_463 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_462 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_461 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_29 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_116 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_115 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_114 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_113 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_929 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_930 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_465 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_930 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_929 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_931 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_932 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_466 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_932 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_931 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_933 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_934 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_467 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_934 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_933 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_935 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_936 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_468 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_936 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_935 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_117 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_468 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_467 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_466 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_465 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_937 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_938 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_469 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_938 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_937 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_939 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_940 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_470 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_940 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_939 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_941 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_942 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_471 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_942 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_941 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_943 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_944 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_472 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_944 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_943 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_118 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_472 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_471 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_470 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_469 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_945 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_946 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_473 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_946 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_945 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_947 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_948 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_474 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_948 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_947 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_949 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_950 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_475 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_950 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_949 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_951 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_952 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_476 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_952 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_951 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_119 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_476 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_475 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_474 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_473 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_953 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_954 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_477 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_954 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_953 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_955 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_956 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_478 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_956 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_955 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_957 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_958 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_479 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_958 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_957 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_959 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_960 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_480 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_960 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_959 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_120 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_480 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_479 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_478 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_477 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_30 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_120 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_119 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_118 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_117 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_961 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_962 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_481 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_962 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_961 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_963 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_964 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_482 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_964 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_963 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_965 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_966 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_483 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_966 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_965 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_967 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_968 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_484 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_968 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_967 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_121 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_484 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_483 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_482 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_481 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_969 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_970 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_485 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_970 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_969 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_971 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_972 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_486 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_972 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_971 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_973 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_974 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_487 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_974 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_973 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_975 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_976 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_488 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_976 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_975 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_122 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_488 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_487 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_486 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_485 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_977 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_978 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_489 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_978 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_977 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_979 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_980 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_490 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_980 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_979 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_981 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_982 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_491 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_982 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_981 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_983 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_984 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_492 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_984 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_983 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_123 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_492 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_491 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_490 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_489 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_985 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_986 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_493 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_986 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_985 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_987 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_988 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_494 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_988 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_987 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_989 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_990 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_495 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_990 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_989 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_991 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_992 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_496 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_992 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_991 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_124 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_496 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_495 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_494 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_493 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_31 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_124 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_123 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_122 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_121 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_993 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_994 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_497 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_994 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_993 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_995 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_996 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_498 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_996 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_995 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_997 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_998 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_499 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_998 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_997 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_999 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1000 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_500 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1000 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_999 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_125 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_500 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_499 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_498 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_497 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1001 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1002 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_501 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1002 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1001 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1003 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1004 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_502 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1004 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1003 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1005 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1006 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_503 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1006 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1005 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1007 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1008 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_504 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1008 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1007 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_126 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_504 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_503 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_502 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_501 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1009 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1010 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_505 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1010 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1009 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1011 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1012 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_506 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1012 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1011 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1013 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1014 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_507 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1014 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1013 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1015 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1016 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_508 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1016 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1015 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_127 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_508 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_507 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_506 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_505 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1017 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1018 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_509 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1018 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1017 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1019 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1020 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_510 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1020 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1019 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1021 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1022 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_511 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1022 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1021 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1023 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1024 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_512 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1024 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1023 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_128 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_512 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_511 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_510 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_509 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_32 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_128 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_127 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_126 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_125 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_8 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n4, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_32 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_31 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_30 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_29 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in8), .Z(n4) );
  CAOR2X1 U6 ( .A(s84[3]), .B(n5), .C(s83[3]), .D(n1), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n5), .C(s83[2]), .D(n1), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n5), .C(s83[1]), .D(n1), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n5), .C(s83[0]), .D(n1), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n4), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n4), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n4), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n4), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n5), .C(c_out810), .D(n1), .Z(c_out8) );
  CANR2X1 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n4), .Z(n1) );
endmodule


module bit32_2 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   c1, c2, c3, n1, n2, n3, n4, n5;

  bit8_8 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8(a32[7:0]), .b8(b32[7:0]), 
        .c_in8(c_in32) );
  bit8_7 A322 ( .sum8(sum32[15:8]), .c_out8(c2), .a8({a32[15:12], n1, 
        a32[10:8]}), .b8(b32[15:8]), .c_in8(c1) );
  bit8_6 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8({a32[23:21], n5, 
        a32[19:16]}), .b8(b32[23:16]), .c_in8(c2) );
  bit8_5 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8({a32[31:27], n3, 
        a32[25:24]}), .b8(b32[31:24]), .c_in8(c3) );
  CNIVX4 U1 ( .A(a32[11]), .Z(n1) );
  CIVX1 U2 ( .A(a32[26]), .Z(n2) );
  CIVX4 U3 ( .A(n2), .Z(n3) );
  CIVX2 U4 ( .A(a32[20]), .Z(n4) );
  CIVX4 U5 ( .A(n4), .Z(n5) );
endmodule


module Add_half_1025 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1026 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_513 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1026 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1025 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1027 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1028 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_514 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1028 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1027 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1029 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1030 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_515 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1030 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1029 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1031 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1032 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_516 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1032 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1031 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_129 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_516 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_515 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_514 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_513 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CIVX1 U5 ( .A(n2), .Z(n3) );
  CMX2XL U6 ( .A0(c_out10), .A1(c_out11), .S(n3), .Z(c_out2) );
  CMX2X1 U7 ( .A0(s3), .A1(s4), .S(n3), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_1033 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1034 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_517 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1034 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1033 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1035 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1036 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_518 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1036 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1035 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1037 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1038 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_519 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1038 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1037 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1039 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1040 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_520 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1040 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1039 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_130 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_520 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_519 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_518 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_517 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(s1), .Z(n3) );
  CIVX2 U8 ( .A(s2), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_1041 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1042 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_521 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1042 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1041 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1043 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1044 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_522 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1044 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1043 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1045 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1046 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_523 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1046 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1045 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1047 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1048 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_524 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1048 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1047 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_131 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_524 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_523 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_522 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_521 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMXI2XL U4 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module Add_half_1049 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1050 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_525 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1050 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1049 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1051 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1052 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_526 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1052 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1051 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1053 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1054 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_527 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1054 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1053 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1055 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1056 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_528 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1056 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1055 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_132 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_528 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_527 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_526 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_525 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMXI2X1 U6 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U7 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module bit4_33 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_132 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_131 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_130 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_129 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CND2X1 U3 ( .A(s44[0]), .B(n5), .Z(n3) );
  CND2X1 U4 ( .A(n2), .B(n3), .Z(sum4[2]) );
  CND2X1 U5 ( .A(s43[0]), .B(n1), .Z(n2) );
  CIVXL U6 ( .A(n5), .Z(n1) );
  CNIVXL U7 ( .A(n5), .Z(n4) );
  CMX2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n5) );
  CIVX1 U9 ( .A(s41[0]), .Z(n7) );
  CIVX1 U10 ( .A(s44[1]), .Z(n8) );
  CIVX1 U11 ( .A(s43[1]), .Z(n9) );
  CMX2XL U12 ( .A0(c_out410), .A1(c_out411), .S(n4), .Z(c_out4) );
  CMX2X1 U13 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U14 ( .A(s42[0]), .Z(n6) );
  CMXI2X1 U15 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[0]) );
  CMXI2X1 U16 ( .A0(n9), .A1(n8), .S(n4), .Z(sum4[3]) );
endmodule


module Add_half_1057 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1058 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_529 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1058 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1057 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1059 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1060 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_530 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1060 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1059 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1061 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1062 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_531 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1062 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1061 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1063 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1064 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_532 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1064 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1063 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_133 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_532 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_531 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_530 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_529 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2XL U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s3), .Z(n4) );
  CIVX2 U9 ( .A(s4), .Z(n3) );
endmodule


module Add_half_1065 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n1) );
  CENX1 U3 ( .A(a), .B(n1), .Z(sum) );
endmodule


module Add_half_1066 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_533 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1066 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1065 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1067 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1068 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_534 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1068 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1067 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1069 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1070 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_535 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1070 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1069 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1071 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1072 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_536 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1072 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1071 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_134 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_536 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_535 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_534 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_533 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_1073 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1074 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_537 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1074 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1073 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1075 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1076 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_538 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1076 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1075 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1077 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1078 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_539 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1078 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1077 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1079 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1080 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVXL U1 ( .A(a), .Z(n1) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_540 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1080 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1079 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_135 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_540 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_539 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_538 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_537 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U4 ( .A(n1), .Z(n4) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_1081 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1082 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_541 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1082 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1081 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1083 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1084 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVX1 U1 ( .A(a), .Z(n1) );
  CND2XL U2 ( .A(n1), .B(b), .Z(n4) );
  CIVXL U3 ( .A(b), .Z(n2) );
  CND2XL U4 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U5 ( .A(n3), .B(n4), .Z(sum) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_542 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1084 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1083 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1085 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1086 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVXL U1 ( .A(a), .Z(n1) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CND2XL U3 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_543 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1086 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1085 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1087 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1088 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVX1 U1 ( .A(b), .Z(n2) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(a), .Z(n1) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_544 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1088 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1087 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_136 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_544 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_543 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_542 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_541 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CIVX1 U5 ( .A(n2), .Z(n7) );
  CIVX1 U6 ( .A(s1), .Z(n6) );
  CMXI2X1 U7 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CMX2XL U8 ( .A0(s3), .A1(s4), .S(n7), .Z(sum2[1]) );
  CIVX2 U9 ( .A(c_out10), .Z(n4) );
  CIVX2 U10 ( .A(c_out11), .Z(n3) );
  CIVX2 U11 ( .A(s2), .Z(n5) );
  CMXI2X1 U12 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
endmodule


module bit4_34 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_136 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_135 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_134 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_133 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMX2X1 U4 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CIVX1 U5 ( .A(s41[1]), .Z(n3) );
  CMX2XL U6 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CMX2X1 U7 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U8 ( .A(s42[1]), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U10 ( .A(s43[0]), .Z(n5) );
  CIVX2 U11 ( .A(s44[0]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(n1), .Z(sum4[2]) );
endmodule


module Add_half_1089 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1090 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_545 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1090 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1089 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1091 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1092 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX2 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_546 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1092 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1091 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1093 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1094 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_547 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1094 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1093 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_1095 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1096 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_548 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1096 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1095 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_137 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_548 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_547 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_546 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_545 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CIVXL U4 ( .A(n2), .Z(n3) );
  CMX2X1 U5 ( .A0(c_out11), .A1(c_out10), .S(n2), .Z(c_out2) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n3), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_1097 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1098 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_549 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1098 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1097 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1099 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1100 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_550 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1100 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1099 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1101 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1102 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2, n3, n4, n5;

  CIVDXL U1 ( .A(b), .Z0(n3) );
  CIVX1 U2 ( .A(a), .Z(n2) );
  CND2X1 U3 ( .A(a), .B(n3), .Z(n4) );
  CND2XL U4 ( .A(n2), .B(b), .Z(n5) );
  CND2X1 U5 ( .A(n4), .B(n5), .Z(sum) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_551 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1102 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1101 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CND2X1 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_1103 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX2 U2 ( .A(n2), .B(b), .Z(sum) );
  CIVXL U3 ( .A(a), .Z(n1) );
  CIVX1 U4 ( .A(n1), .Z(n2) );
endmodule


module Add_half_1104 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2, n3, n4, n5;

  CND2XL U1 ( .A(n2), .B(b), .Z(n5) );
  CIVDXL U2 ( .A(b), .Z0(n3) );
  CND2X1 U3 ( .A(a), .B(n3), .Z(n4) );
  CIVX1 U4 ( .A(a), .Z(n2) );
  CND2X1 U5 ( .A(n4), .B(n5), .Z(sum) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_552 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1104 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1103 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_138 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_552 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_551 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_550 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_549 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n3) );
  CMX2X1 U4 ( .A0(c_out11), .A1(c_out10), .S(n1), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out01), .A1(c_out00), .S(n3), .Z(n1) );
  CMX2XL U6 ( .A0(c_out01), .A1(c_out00), .S(n3), .Z(n2) );
  CIVX1 U7 ( .A(s2), .Z(n4) );
  CMXI2X1 U8 ( .A0(n7), .A1(n6), .S(n2), .Z(sum2[1]) );
  CIVX1 U9 ( .A(s3), .Z(n7) );
  CIVX2 U10 ( .A(s1), .Z(n5) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
endmodule


module Add_half_1105 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1106 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_553 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1106 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1105 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1107 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1108 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_554 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1108 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1107 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1109 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CEOXL U2 ( .A(b), .B(n1), .Z(sum) );
  CND2X2 U3 ( .A(a), .B(b), .Z(n2) );
  CIVX2 U4 ( .A(n2), .Z(c_out) );
endmodule


module Add_half_1110 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_555 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1110 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1109 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_1111 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CND2X2 U2 ( .A(a), .B(b), .Z(n2) );
  CEOXL U3 ( .A(b), .B(n1), .Z(sum) );
  CIVX2 U4 ( .A(n2), .Z(c_out) );
endmodule


module Add_half_1112 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_556 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1112 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1111 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_139 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8, n9;

  Add_full_556 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_555 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_554 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_553 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CIVX1 U4 ( .A(s4), .Z(n8) );
  CIVX1 U5 ( .A(s3), .Z(n9) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n3) );
  CMX2XL U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMXI2X1 U8 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CIVX1 U9 ( .A(s2), .Z(n6) );
  CIVX1 U10 ( .A(s1), .Z(n7) );
  CMXI2XL U11 ( .A0(n9), .A1(n8), .S(n2), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_out10), .Z(n5) );
  CIVX2 U13 ( .A(c_out11), .Z(n4) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_1113 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1114 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_557 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1114 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1113 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1115 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1116 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_558 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1116 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1115 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1117 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3;

  CENX1 U1 ( .A(n1), .B(n3), .Z(sum) );
  CIVX2 U2 ( .A(n2), .Z(c_out) );
  CND2X2 U3 ( .A(a), .B(b), .Z(n2) );
  CNIVXL U4 ( .A(a), .Z(n1) );
  CIVX2 U5 ( .A(b), .Z(n3) );
endmodule


module Add_half_1118 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_559 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1118 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1117 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_1119 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVX2 U1 ( .A(b), .Z(n3) );
  CIVXL U2 ( .A(a), .Z(n1) );
  CIVXL U3 ( .A(n1), .Z(n2) );
  CND2IX2 U4 ( .B(n3), .A(a), .Z(n4) );
  CEOXL U5 ( .A(b), .B(n2), .Z(sum) );
  CIVX2 U6 ( .A(n4), .Z(c_out) );
endmodule


module Add_half_1120 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_560 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1120 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1119 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_140 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_560 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_559 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_558 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_557 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s4), .Z(n5) );
  CIVX1 U4 ( .A(s3), .Z(n6) );
  CMX2XL U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U6 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMX2XL U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2XL U8 ( .A0(n6), .A1(n5), .S(n1), .Z(sum2[1]) );
  CIVX2 U9 ( .A(c_out10), .Z(n4) );
  CIVX2 U10 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U11 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module bit4_35 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_140 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_139 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_138 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_137 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(n4), .Z(n1) );
  CIVXL U4 ( .A(n4), .Z(n9) );
  CIVX1 U5 ( .A(c_out410), .Z(n6) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n4) );
  CIVXL U7 ( .A(n9), .Z(n2) );
  CIVX1 U8 ( .A(n2), .Z(n3) );
  CIVX1 U9 ( .A(c_out411), .Z(n5) );
  CMXI2X1 U10 ( .A0(n6), .A1(n5), .S(n1), .Z(c_out4) );
  CMX2X1 U11 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U12 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMXI2XL U13 ( .A0(n11), .A1(n10), .S(n3), .Z(sum4[3]) );
  CMXI2XL U14 ( .A0(n8), .A1(n7), .S(n9), .Z(sum4[2]) );
  CIVX2 U15 ( .A(s43[0]), .Z(n8) );
  CIVX2 U16 ( .A(s44[0]), .Z(n7) );
  CIVX2 U17 ( .A(s43[1]), .Z(n11) );
  CIVX2 U18 ( .A(s44[1]), .Z(n10) );
endmodule


module Add_half_1121 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1122 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_561 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1122 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1121 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1123 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1124 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_562 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1124 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1123 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1125 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1126 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_563 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1126 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1125 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1127 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1128 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_564 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1128 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1127 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_141 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_564 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_563 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_562 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_561 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n3) );
  CMX2XL U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMX2X1 U6 ( .A0(c_out11), .A1(c_out10), .S(n3), .Z(c_out2) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(s3), .Z(n5) );
  CIVX2 U9 ( .A(s4), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_1129 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1130 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_565 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1130 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1129 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1131 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1132 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_566 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1132 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1131 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1133 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1134 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(a), .B(n2), .Z(n3) );
  CND2XL U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_567 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1134 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1133 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1135 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1136 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_568 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1136 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1135 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_142 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_568 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_567 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_566 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_565 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n2) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n3) );
  CMX2XL U5 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CMX2X1 U6 ( .A0(c_out11), .A1(c_out10), .S(n3), .Z(c_out2) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(s3), .Z(n5) );
  CIVX2 U9 ( .A(s4), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
endmodule


module Add_half_1137 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1138 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_569 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1138 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1137 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1139 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1140 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_570 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1140 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1139 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1141 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1142 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_571 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1142 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1141 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_1143 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1144 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_572 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1144 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1143 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_143 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_572 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_571 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_570 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_569 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX1 U4 ( .A(c_out11), .Z(n2) );
  CIVX2 U5 ( .A(n1), .Z(n4) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_1145 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1146 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_573 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1146 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1145 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1147 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1148 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_574 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1148 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1147 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1149 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1150 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_575 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1150 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1149 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_1151 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1152 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_576 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1152 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1151 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_144 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_576 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_575 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_574 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_573 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s4), .Z(n5) );
  CIVX1 U4 ( .A(s3), .Z(n6) );
  CIVX2 U5 ( .A(n1), .Z(n4) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2XL U7 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U8 ( .A(c_out10), .Z(n3) );
  CIVX2 U9 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U10 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_36 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_144 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_143 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_142 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_141 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CIVX2 U4 ( .A(c_in4), .Z(n1) );
  CIVX1 U5 ( .A(c_out411), .Z(n4) );
  CMXI2X1 U6 ( .A0(c_out401), .A1(c_out400), .S(n1), .Z(n3) );
  CMXI2X1 U7 ( .A0(n11), .A1(n10), .S(n2), .Z(sum4[2]) );
  CIVX1 U8 ( .A(s41[1]), .Z(n9) );
  CIVX1 U9 ( .A(s43[0]), .Z(n11) );
  CMXI2X1 U10 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out4) );
  CIVX2 U11 ( .A(c_out410), .Z(n5) );
  CMXI2XL U12 ( .A0(n13), .A1(n12), .S(n2), .Z(sum4[3]) );
  CIVX2 U13 ( .A(s41[0]), .Z(n7) );
  CIVX2 U14 ( .A(s42[0]), .Z(n6) );
  CMXI2X1 U15 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U16 ( .A(s42[1]), .Z(n8) );
  CMXI2X1 U17 ( .A0(n9), .A1(n8), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U18 ( .A(s44[0]), .Z(n10) );
  CIVX2 U19 ( .A(s43[1]), .Z(n13) );
  CIVX2 U20 ( .A(s44[1]), .Z(n12) );
endmodule


module bit8_9 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, net68843, net85358, net89638,
         net90064, net95571, net97521, net111077, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_36 A81 ( .sum4(s81), .c_out4(c_out800), .a4({a8[3:1], n22}), .b4({n1, 
        b8[2:0]}), .c_in4(1'b0) );
  bit4_35 A82 ( .sum4(s82), .c_out4(c_out801), .a4({a8[3:1], n8}), .b4({n1, 
        b8[2:0]}), .c_in4(1'b1) );
  bit4_34 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4({n21, b8[6:4]}), .c_in4(1'b0) );
  bit4_33 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4({n21, b8[6:4]}), .c_in4(1'b1) );
  CIVX3 U3 ( .A(n4), .Z(sum8[6]) );
  CIVX1 U4 ( .A(net68843), .Z(net95571) );
  CIVX2 U5 ( .A(net90064), .Z(net97521) );
  CNIVX4 U6 ( .A(b8[3]), .Z(n1) );
  CND2X1 U7 ( .A(s81[1]), .B(net111077), .Z(n2) );
  CND2X1 U8 ( .A(s82[1]), .B(net85358), .Z(n3) );
  CND2X2 U9 ( .A(n2), .B(n3), .Z(sum8[1]) );
  CND2X1 U10 ( .A(s81[2]), .B(net111077), .Z(n6) );
  CIVX2 U11 ( .A(n10), .Z(n14) );
  CNIVX1 U12 ( .A(n18), .Z(n9) );
  CMXI2X1 U13 ( .A0(s84[2]), .A1(s83[2]), .S(n18), .Z(n4) );
  CMX2X1 U14 ( .A0(s82[0]), .A1(s81[0]), .S(n5), .Z(sum8[0]) );
  CIVX2 U15 ( .A(c_in8), .Z(n5) );
  CIVX2 U16 ( .A(n5), .Z(net90064) );
  CIVX2 U17 ( .A(n5), .Z(net85358) );
  CND2X4 U18 ( .A(n12), .B(n13), .Z(sum8[5]) );
  CND2XL U19 ( .A(s82[2]), .B(net85358), .Z(n7) );
  CND2X2 U20 ( .A(n7), .B(n6), .Z(sum8[2]) );
  CIVX1 U21 ( .A(net85358), .Z(net111077) );
  CMX2X2 U22 ( .A0(s84[3]), .A1(s83[3]), .S(n9), .Z(sum8[7]) );
  CNIVX4 U23 ( .A(a8[0]), .Z(n8) );
  CND2X2 U24 ( .A(n25), .B(s83[0]), .Z(n16) );
  CANR2X1 U25 ( .A(net97521), .B(c_out800), .C(net85358), .D(c_out801), .Z(n10) );
  CND2X2 U26 ( .A(n11), .B(s84[1]), .Z(n12) );
  CND2X1 U27 ( .A(s83[1]), .B(n17), .Z(n13) );
  CIVX1 U28 ( .A(n17), .Z(n11) );
  CND2X4 U29 ( .A(n15), .B(n16), .Z(sum8[4]) );
  CND2X2 U30 ( .A(n14), .B(s84[0]), .Z(n15) );
  CANR2X1 U31 ( .A(c_out800), .B(net68843), .C(net85358), .D(c_out801), .Z(n25) );
  CANR2X1 U32 ( .A(net97521), .B(c_out800), .C(c_out801), .D(net95571), .Z(n17) );
  CANR2X1 U33 ( .A(net97521), .B(c_out800), .C(net85358), .D(c_out801), .Z(n18) );
  CND2XL U34 ( .A(s82[3]), .B(net95571), .Z(n20) );
  CND2X1 U35 ( .A(s81[3]), .B(net89638), .Z(n19) );
  CND2X2 U36 ( .A(n19), .B(n20), .Z(sum8[3]) );
  CIVXL U37 ( .A(net95571), .Z(net89638) );
  CNIVX4 U38 ( .A(b8[7]), .Z(n21) );
  CNIVX4 U39 ( .A(a8[0]), .Z(n22) );
  CMXI2XL U40 ( .A0(n24), .A1(n23), .S(n9), .Z(c_out8) );
  CIVX2 U41 ( .A(c_out811), .Z(n24) );
  CIVX2 U42 ( .A(c_out810), .Z(n23) );
  CIVX2 U43 ( .A(net90064), .Z(net68843) );
endmodule


module Add_half_1153 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1154 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_577 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1154 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1153 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1155 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1156 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_578 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1156 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1155 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1157 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOX1 U1 ( .A(b), .B(n1), .Z(sum) );
  CNIVXL U2 ( .A(a), .Z(n1) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1158 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CENX1 U1 ( .A(n1), .B(b), .Z(sum) );
  CIVX1 U2 ( .A(a), .Z(n1) );
  CIVXL U3 ( .A(n1), .Z(n2) );
  CAN2XL U4 ( .A(b), .B(n2), .Z(c_out) );
endmodule


module Add_full_579 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1158 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1157 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1159 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOX1 U1 ( .A(b), .B(n1), .Z(sum) );
  CNIVXL U2 ( .A(a), .Z(n1) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1160 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_580 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1160 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1159 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_145 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_580 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_579 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_578 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_577 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2X1 U3 ( .A(c_out11), .B(n1), .Z(n2) );
  CND2X1 U4 ( .A(c_out10), .B(n6), .Z(n3) );
  CND2X2 U5 ( .A(n2), .B(n3), .Z(c_out2) );
  CIVX2 U6 ( .A(n6), .Z(n1) );
  CIVX2 U7 ( .A(c_in2), .Z(n4) );
  CMX2XL U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U9 ( .A0(c_out01), .A1(c_out00), .S(n4), .Z(n6) );
  CMX2XL U10 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n5) );
  CMXI2XL U11 ( .A0(n8), .A1(n7), .S(n5), .Z(sum2[1]) );
  CIVX2 U12 ( .A(s3), .Z(n8) );
  CIVX2 U13 ( .A(s4), .Z(n7) );
endmodule


module Add_half_1161 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1162 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENXL U1 ( .A(a), .B(b), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_581 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1162 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1161 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1163 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1164 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_582 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1164 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1163 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1165 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(n1), .Z(sum) );
endmodule


module Add_half_1166 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_583 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1166 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1165 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_1167 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(b), .B(n1), .Z(sum) );
  CNIVXL U2 ( .A(a), .Z(n1) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1168 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_584 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1168 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1167 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_146 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_584 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_583 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_582 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_581 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMX2X1 U5 ( .A0(c_out11), .A1(c_out10), .S(n2), .Z(c_out2) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module Add_half_1169 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1170 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_585 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1170 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1169 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1171 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1172 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_586 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1172 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1171 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1173 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3;

  CIVX2 U1 ( .A(a), .Z(n2) );
  CNR2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n1) );
  CIVX1 U4 ( .A(n2), .Z(n3) );
  CEOXL U5 ( .A(b), .B(n3), .Z(sum) );
endmodule


module Add_half_1174 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVXL U1 ( .A(b), .Z(n2) );
  CIVX1 U2 ( .A(a), .Z(n1) );
  CND2X1 U3 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CND2XL U5 ( .A(a), .B(n2), .Z(n3) );
  CAN2XL U6 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_587 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1174 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1173 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1175 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1176 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_588 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1176 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1175 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_147 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_588 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_587 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_586 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_585 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(c_out11), .Z(n3) );
  CMX2XL U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U5 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out10), .Z(n4) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module Add_half_1177 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1178 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_589 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1178 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1177 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1179 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1180 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_590 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1180 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1179 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1181 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(n2) );
  CEOXL U3 ( .A(b), .B(n2), .Z(sum) );
  CAN2X1 U4 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1182 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n1), .B(b), .Z(n4) );
  CIVX1 U2 ( .A(b), .Z(n2) );
  CIVX1 U3 ( .A(a), .Z(n1) );
  CND2XL U4 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U5 ( .A(n4), .B(n3), .Z(sum) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_591 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1182 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1181 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1183 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(n2) );
  CEOXL U3 ( .A(b), .B(n2), .Z(sum) );
  CAN2X1 U4 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1184 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U2 ( .A(n4), .B(n3), .Z(sum) );
  CND2XL U3 ( .A(a), .B(n2), .Z(n3) );
  CIVX1 U4 ( .A(b), .Z(n2) );
  CIVX1 U5 ( .A(a), .Z(n1) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_592 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1184 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1183 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_148 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_592 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_591 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_590 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_589 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n7), .A1(n6), .S(n1), .Z(c_out2) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CNIVXL U5 ( .A(c_out00), .Z(n2) );
  CIVX2 U6 ( .A(c_in2), .Z(n5) );
  CMX2X1 U7 ( .A0(n4), .A1(n2), .S(n5), .Z(n3) );
  CIVX1 U8 ( .A(c_out10), .Z(n7) );
  CIVX1 U9 ( .A(c_out11), .Z(n6) );
  CMX2X1 U10 ( .A0(s3), .A1(s4), .S(n3), .Z(sum2[1]) );
  CNIVXL U11 ( .A(c_out01), .Z(n4) );
  CMX2X1 U12 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module bit4_37 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_148 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_147 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_146 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_145 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CND2X2 U3 ( .A(n2), .B(n3), .Z(n1) );
  CND2X2 U4 ( .A(c_out401), .B(c_in4), .Z(n2) );
  CND2X2 U5 ( .A(n3), .B(n2), .Z(n4) );
  CMX2X1 U6 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CND2X2 U7 ( .A(c_out400), .B(n5), .Z(n3) );
  CIVXL U8 ( .A(s44[0]), .Z(n11) );
  CIVXL U9 ( .A(s43[0]), .Z(n12) );
  CMXI2XL U10 ( .A0(n12), .A1(n11), .S(n1), .Z(sum4[2]) );
  CIVX2 U11 ( .A(n1), .Z(n6) );
  CIVX2 U12 ( .A(c_in4), .Z(n5) );
  CND2X2 U13 ( .A(c_out411), .B(n4), .Z(n8) );
  CND2X2 U14 ( .A(c_out410), .B(n6), .Z(n7) );
  CND2X2 U15 ( .A(n7), .B(n8), .Z(c_out4) );
  CMX2X1 U16 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U17 ( .A(s41[0]), .Z(n10) );
  CIVX2 U18 ( .A(s42[0]), .Z(n9) );
  CMXI2X1 U19 ( .A0(n10), .A1(n9), .S(c_in4), .Z(sum4[0]) );
endmodule


module Add_half_1185 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1186 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENXL U1 ( .A(a), .B(b), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_593 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1186 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1185 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1187 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1188 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_594 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1188 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1187 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1189 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1190 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_595 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1190 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1189 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_1191 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1192 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_596 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1192 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1191 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_149 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_596 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_595 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_594 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_593 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CIVX2 U5 ( .A(n2), .Z(n5) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(c_out10), .A1(c_out11), .S(n5), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n4) );
  CIVX2 U9 ( .A(s2), .Z(n3) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_1193 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1194 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_597 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1194 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1193 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1195 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1196 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_598 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1196 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1195 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1197 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n4;

  CENX1 U1 ( .A(n2), .B(n4), .Z(sum) );
  CIVXL U2 ( .A(a), .Z(n1) );
  CIVXL U3 ( .A(n1), .Z(n2) );
  CAN2X1 U4 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U5 ( .A(b), .Z(n4) );
endmodule


module Add_half_1198 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n1), .B(b), .Z(n4) );
  CIVXL U2 ( .A(a), .Z(n1) );
  CIVXL U3 ( .A(b), .Z(n2) );
  CND2XL U4 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U5 ( .A(n3), .B(n4), .Z(sum) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_599 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1198 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1197 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_1199 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1200 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_600 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1200 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1199 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_150 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_600 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_599 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_598 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_597 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2XL U3 ( .A(c_out10), .B(n3), .Z(n1) );
  CND2XL U4 ( .A(n4), .B(c_out11), .Z(n2) );
  CND2X1 U5 ( .A(n1), .B(n2), .Z(c_out2) );
  CIVX1 U6 ( .A(n3), .Z(n4) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CMX2XL U8 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U9 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_1201 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1202 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_601 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1202 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1201 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1203 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1204 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_602 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1204 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1203 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1205 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1206 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_603 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1206 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1205 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1207 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(n2) );
  CEOXL U3 ( .A(b), .B(n2), .Z(sum) );
  CAN2X1 U4 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1208 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n4), .B(n3), .Z(sum) );
  CND2X1 U3 ( .A(n1), .B(b), .Z(n4) );
  CIVXL U4 ( .A(b), .Z(n2) );
  CIVX1 U5 ( .A(a), .Z(n1) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_604 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1208 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1207 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_151 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_604 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_603 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_602 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_601 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n2) );
  CMX2XL U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U5 ( .A(c_out10), .Z(n5) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n3) );
  CIVX1 U7 ( .A(c_out11), .Z(n4) );
  CIVX1 U8 ( .A(s2), .Z(n6) );
  CIVX1 U9 ( .A(s1), .Z(n7) );
  CMXI2X1 U10 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CMX2XL U11 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMXI2X1 U12 ( .A0(n7), .A1(n6), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_1209 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1210 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_605 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1210 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1209 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1211 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1212 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_606 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1212 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1211 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1213 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1214 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_607 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1214 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1213 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1215 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CEOXL U2 ( .A(b), .B(n1), .Z(sum) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1216 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_608 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1216 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1215 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_152 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_608 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_607 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_606 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_605 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(c_out10), .Z(n4) );
  CIVX1 U4 ( .A(s3), .Z(n6) );
  CIVX1 U5 ( .A(c_out11), .Z(n3) );
  CMX2XL U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U7 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2XL U9 ( .A0(n6), .A1(n5), .S(n1), .Z(sum2[1]) );
  CMXI2X1 U10 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module bit4_38 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_152 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_151 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_150 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_149 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CND2IX1 U3 ( .B(n3), .A(c_out411), .Z(n1) );
  CMX2X2 U4 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n4) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n3) );
  CND2X1 U6 ( .A(n3), .B(c_out410), .Z(n2) );
  CND2X2 U7 ( .A(n1), .B(n2), .Z(c_out4) );
  CMX2X1 U8 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2XL U9 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2X1 U10 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U11 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
endmodule


module Add_half_1217 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1218 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_609 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1218 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1217 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1219 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1220 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_610 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1220 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1219 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1221 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CEOXL U3 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1222 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_611 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1222 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1221 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1223 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CEOXL U3 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1224 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_612 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1224 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1223 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_153 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_612 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_611 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_610 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_609 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n4) );
  CMXI2XL U4 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module Add_half_1225 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CENX1 U4 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1226 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_613 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1226 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1225 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1227 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1228 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_614 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1228 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1227 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1229 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CNIVX1 U1 ( .A(a), .Z(n1) );
  CIVX1 U2 ( .A(n2), .Z(c_out) );
  CEOXL U3 ( .A(n1), .B(b), .Z(sum) );
  CND2X1 U4 ( .A(a), .B(b), .Z(n2) );
endmodule


module Add_half_1230 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n1), .B(b), .Z(n4) );
  CIVX2 U2 ( .A(a), .Z(n1) );
  CND2XL U3 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_615 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1230 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1229 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1231 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1232 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_616 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1232 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1231 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_154 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_616 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_615 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_614 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_613 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_1233 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1234 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_617 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1234 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1233 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1235 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1236 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_618 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1236 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1235 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1237 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1238 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVX1 U1 ( .A(a), .Z(n1) );
  CND2X1 U2 ( .A(n1), .B(b), .Z(n4) );
  CIVX1 U3 ( .A(b), .Z(n2) );
  CND2X1 U4 ( .A(a), .B(n2), .Z(n3) );
  CND2X2 U5 ( .A(n3), .B(n4), .Z(sum) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_619 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1238 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1237 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1239 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1240 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_620 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1240 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1239 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_155 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n2, n3, n4, n5;

  Add_full_620 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_619 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_618 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_617 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CIVDXL U4 ( .A(n2), .Z0(n5) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n4) );
  CIVX2 U8 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module Add_half_1241 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1242 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_621 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1242 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1241 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1243 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1244 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_622 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1244 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1243 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1245 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1246 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_623 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1246 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1245 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1247 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1248 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n3), .B(n4), .Z(sum) );
  CND2X1 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2XL U3 ( .A(a), .B(n2), .Z(n3) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_624 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1248 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1247 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_156 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_624 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_623 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_622 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_621 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n2) );
  CMX2XL U4 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CMXI2X1 U5 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n3) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CIVX2 U8 ( .A(c_out10), .Z(n5) );
  CIVX2 U9 ( .A(c_out11), .Z(n4) );
  CIVX2 U10 ( .A(s1), .Z(n7) );
  CIVX2 U11 ( .A(s2), .Z(n6) );
  CMXI2X1 U12 ( .A0(n7), .A1(n6), .S(c_in2), .Z(sum2[0]) );
endmodule


module bit4_39 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_156 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_155 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_154 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_153 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX1 U4 ( .A(c_out410), .Z(n4) );
  CIVX1 U5 ( .A(c_out411), .Z(n3) );
  CMXI2X1 U6 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out4) );
  CMX2XL U7 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U8 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U9 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMXI2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CIVX2 U11 ( .A(s43[0]), .Z(n6) );
  CIVX2 U12 ( .A(s44[0]), .Z(n5) );
  CMXI2X1 U13 ( .A0(n6), .A1(n5), .S(n1), .Z(sum4[2]) );
endmodule


module Add_half_1249 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1250 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_625 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1250 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1249 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1251 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1252 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_626 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1252 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1251 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1253 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1254 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_627 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1254 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1253 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1255 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1256 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_628 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1256 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1255 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_157 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_628 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_627 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_626 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_625 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n6) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_1257 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1258 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_629 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1258 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1257 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1259 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1260 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_630 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1260 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1259 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1261 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1262 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_631 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1262 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1261 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1263 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1264 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_632 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1264 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1263 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_158 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_632 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_631 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_630 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_629 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CIVX1 U4 ( .A(n2), .Z(n5) );
  CMXI2X1 U5 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out10), .Z(n4) );
  CIVX2 U9 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(n5), .Z(c_out2) );
endmodule


module Add_half_1265 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CENX1 U4 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1266 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_633 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1266 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1265 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_1267 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1268 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_634 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1268 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1267 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1269 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net89574;
  assign c_out = net89574;

  CAN2X1 U1 ( .A(b), .B(a), .Z(net89574) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1270 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88859;
  assign c_out = net88859;

  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(net88859) );
endmodule


module Add_full_635 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1270 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1269 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n1), .B(n2), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n2) );
  CIVX2 U3 ( .A(w3), .Z(n1) );
endmodule


module Add_half_1271 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CND2X1 U2 ( .A(b), .B(a), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1272 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_636 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1272 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1271 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_159 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, net113874,
         net113873, net69310, n1, n2, n3;

  Add_full_636 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_635 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_634 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_633 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s3), .A1(s4), .S(net113874), .Z(sum2[1]) );
  CMXI2X1 U4 ( .A0(n1), .A1(n2), .S(net69310), .Z(c_out2) );
  CIVX2 U5 ( .A(n3), .Z(net69310) );
  CIVXL U6 ( .A(net69310), .Z(net113873) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CIVX2 U9 ( .A(c_out10), .Z(n1) );
  CMX2X1 U10 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX1 U11 ( .A(net113873), .Z(net113874) );
endmodule


module Add_half_1273 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1274 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_637 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1274 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1273 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1275 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1276 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_638 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1276 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1275 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1277 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1278 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_639 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1278 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1277 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1279 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1280 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_640 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1280 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1279 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_160 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_640 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_639 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_638 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_637 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n4), .A1(n5), .S(n1), .Z(sum2[1]) );
  CMXI2X1 U4 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
endmodule


module bit4_40 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, net69344, net69345, net69351,
         net69352, net69346, n1, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_160 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_159 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_158 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_157 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2XL U4 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n5) );
  CMX2XL U5 ( .A0(s43[0]), .A1(s44[0]), .S(net69346), .Z(sum4[2]) );
  CND2X2 U6 ( .A(c_out411), .B(net69346), .Z(n4) );
  CND2X2 U7 ( .A(n4), .B(n3), .Z(c_out4) );
  CND2XL U8 ( .A(n5), .B(c_out410), .Z(n3) );
  CIVX2 U9 ( .A(n1), .Z(net69346) );
  CMXI2X1 U10 ( .A0(net69351), .A1(net69352), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U11 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMXI2XL U12 ( .A0(net69344), .A1(net69345), .S(net69346), .Z(sum4[3]) );
  CIVX2 U13 ( .A(s41[0]), .Z(net69351) );
  CIVX2 U14 ( .A(s42[0]), .Z(net69352) );
  CIVX2 U15 ( .A(s43[1]), .Z(net69344) );
  CIVX2 U16 ( .A(s44[1]), .Z(net69345) );
endmodule


module bit8_10 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, net69358, net90529, net92097,
         net99249, net100621, net100615, net102635, net102634, net104733,
         net106308, net95356, net100619, net69374, net69373, net89852, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n24, n25, n26, n27, n28, n29;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;
  assign sum8[1] = net99249;

  bit4_40 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4({b8[3:1], n20}), .c_in4(1'b0) );
  bit4_39 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4({b8[3:1], n20}), .c_in4(1'b1) );
  bit4_38 A83 ( .sum4(s83), .c_out4(c_out810), .a4({a8[7:6], n18, n15}), .b4(
        b8[7:4]), .c_in4(1'b0) );
  bit4_37 A84 ( .sum4(s84), .c_out4(c_out811), .a4({a8[7:6], n16, n22}), .b4(
        b8[7:4]), .c_in4(1'b1) );
  CNIVX3 U3 ( .A(a8[4]), .Z(n15) );
  CND2X2 U4 ( .A(s82[2]), .B(n1), .Z(n2) );
  CND2X1 U5 ( .A(s81[2]), .B(n11), .Z(n3) );
  CND2X4 U6 ( .A(n2), .B(n3), .Z(sum8[2]) );
  CIVX1 U7 ( .A(n11), .Z(n1) );
  CNIVX3 U8 ( .A(a8[4]), .Z(n22) );
  CMXI2X4 U9 ( .A0(n28), .A1(n29), .S(n4), .Z(sum8[7]) );
  CMXI2X1 U10 ( .A0(n26), .A1(n27), .S(n4), .Z(sum8[6]) );
  CIVX3 U11 ( .A(n17), .Z(n16) );
  CND2XL U12 ( .A(net95356), .B(c_out801), .Z(n6) );
  CND2X1 U13 ( .A(n11), .B(c_out800), .Z(n5) );
  CND2X1 U14 ( .A(n5), .B(n6), .Z(n4) );
  CIVX1 U15 ( .A(c_in8), .Z(n7) );
  CIVX1 U16 ( .A(c_in8), .Z(net100619) );
  CIVX1 U17 ( .A(net100621), .Z(net92097) );
  CIVX2 U18 ( .A(n7), .Z(n8) );
  CIVXL U19 ( .A(n11), .Z(n9) );
  CIVXL U20 ( .A(net95356), .Z(n10) );
  CIVX1 U21 ( .A(net100619), .Z(net95356) );
  CIVX2 U22 ( .A(n8), .Z(n11) );
  CMXI2X1 U23 ( .A0(c_out801), .A1(c_out800), .S(n7), .Z(net89852) );
  CMXI2X1 U24 ( .A0(net69373), .A1(net69374), .S(net89852), .Z(c_out8) );
  CANR2X1 U25 ( .A(net92097), .B(c_out800), .C(c_out801), .D(net95356), .Z(
        net69358) );
  CIVXL U26 ( .A(c_out801), .Z(net102634) );
  CNIVXL U27 ( .A(c_out800), .Z(net104733) );
  CIVX2 U28 ( .A(c_out810), .Z(net69374) );
  CIVX2 U29 ( .A(c_out811), .Z(net69373) );
  CIVX3 U30 ( .A(n17), .Z(n18) );
  CMXI2X1 U31 ( .A0(n13), .A1(n14), .S(net100621), .Z(n12) );
  CIVX2 U32 ( .A(n12), .Z(net100615) );
  CNIVX1 U33 ( .A(net95356), .Z(net106308) );
  CMX2X2 U34 ( .A0(s81[1]), .A1(s82[1]), .S(n8), .Z(net99249) );
  CIVX2 U35 ( .A(net100619), .Z(net100621) );
  CIVX2 U36 ( .A(s82[0]), .Z(n14) );
  CIVX2 U37 ( .A(s81[0]), .Z(n13) );
  CIVX3 U38 ( .A(n21), .Z(sum8[5]) );
  CIVX2 U39 ( .A(s83[2]), .Z(n26) );
  CIVX2 U40 ( .A(a8[5]), .Z(n17) );
  CMXI2X1 U41 ( .A0(s84[1]), .A1(s83[1]), .S(net90529), .Z(n21) );
  CIVXL U42 ( .A(net102634), .Z(net102635) );
  CMX2X2 U43 ( .A0(s81[3]), .A1(s82[3]), .S(n9), .Z(sum8[3]) );
  CIVX4 U44 ( .A(net100615), .Z(sum8[0]) );
  CANR2X1 U45 ( .A(net104733), .B(n10), .C(net106308), .D(net102635), .Z(
        net90529) );
  CIVX2 U46 ( .A(b8[0]), .Z(n19) );
  CMXI2X1 U47 ( .A0(n25), .A1(n24), .S(net69358), .Z(sum8[4]) );
  CIVX4 U48 ( .A(n19), .Z(n20) );
  CIVXL U49 ( .A(s84[2]), .Z(n27) );
  CIVX2 U50 ( .A(s84[0]), .Z(n25) );
  CIVX2 U51 ( .A(s83[0]), .Z(n24) );
  CIVX2 U52 ( .A(s84[3]), .Z(n29) );
  CIVX2 U53 ( .A(s83[3]), .Z(n28) );
endmodule


module Add_half_1281 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1282 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_641 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1282 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1281 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1283 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1284 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_642 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1284 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1283 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1285 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1286 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_643 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1286 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1285 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1287 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1288 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_644 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1288 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1287 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_161 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_644 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_643 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_642 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_641 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n4) );
  CMXI2X1 U4 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_1289 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1290 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_645 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1290 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1289 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1291 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1292 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_646 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1292 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1291 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1293 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1294 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_647 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1294 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1293 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1295 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1296 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_648 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1296 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1295 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_162 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_648 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_647 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_646 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_645 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n4), .Z(n3) );
  CND2X1 U4 ( .A(c_out10), .B(n4), .Z(n1) );
  CND2X1 U5 ( .A(c_out11), .B(n3), .Z(n2) );
  CND2X1 U6 ( .A(n1), .B(n2), .Z(c_out2) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n3), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n4) );
endmodule


module Add_half_1297 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1298 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_649 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1298 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1297 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1299 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1300 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_650 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1300 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1299 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1301 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3;

  CIVX2 U1 ( .A(n2), .Z(c_out) );
  CND2IX1 U2 ( .B(n1), .A(a), .Z(n2) );
  CIVX2 U3 ( .A(b), .Z(n1) );
  CNIVXL U4 ( .A(a), .Z(n3) );
  CEOXL U5 ( .A(b), .B(n3), .Z(sum) );
endmodule


module Add_half_1302 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_651 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1302 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1301 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1303 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVX1 U1 ( .A(n2), .Z(c_out) );
  CND2IX1 U2 ( .B(n1), .A(a), .Z(n2) );
  CIVX2 U3 ( .A(b), .Z(n1) );
  CIVXL U4 ( .A(a), .Z(n3) );
  CIVX1 U5 ( .A(n3), .Z(n4) );
  CEOXL U6 ( .A(b), .B(n4), .Z(sum) );
endmodule


module Add_half_1304 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n4), .B(n3), .Z(sum) );
  CIVX1 U2 ( .A(b), .Z(n2) );
  CND2XL U3 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U4 ( .A(n1), .B(b), .Z(n4) );
  CIVXL U5 ( .A(a), .Z(n1) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_652 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1304 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1303 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_163 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8, n9;

  Add_full_652 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_651 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_650 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_649 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(c_out01), .Z(n1) );
  CIVXL U4 ( .A(n1), .Z(n2) );
  CND2X2 U5 ( .A(c_out01), .B(c_in2), .Z(n3) );
  CMX2X1 U6 ( .A0(s3), .A1(s4), .S(n7), .Z(sum2[1]) );
  CMXI2X1 U7 ( .A0(n9), .A1(n8), .S(n5), .Z(c_out2) );
  CND2X2 U8 ( .A(c_out00), .B(n6), .Z(n4) );
  CND2X2 U9 ( .A(n4), .B(n3), .Z(n5) );
  CIVX2 U10 ( .A(c_in2), .Z(n6) );
  CMX2XL U11 ( .A0(c_out00), .A1(n2), .S(c_in2), .Z(n7) );
  CMX2X1 U12 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U13 ( .A(c_out10), .Z(n9) );
  CIVX2 U14 ( .A(c_out11), .Z(n8) );
endmodule


module Add_half_1305 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1306 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_653 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1306 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1305 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1307 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1308 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_654 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1308 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1307 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1309 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVX1 U1 ( .A(a), .Z(n1) );
  CEOXL U2 ( .A(b), .B(n1), .Z(sum) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1310 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X2 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X2 U3 ( .A(n4), .B(n3), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_655 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1310 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1309 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1311 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(n2) );
  CEOXL U3 ( .A(b), .B(n2), .Z(sum) );
  CAN2X1 U4 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1312 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X2 U1 ( .A(n1), .B(b), .Z(n4) );
  CIVX1 U2 ( .A(a), .Z(n1) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
  CND2XL U4 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U5 ( .A(n4), .B(n3), .Z(sum) );
  CIVX1 U6 ( .A(b), .Z(n2) );
endmodule


module Add_full_656 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1312 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1311 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_164 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8, n9;

  Add_full_656 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_655 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_654 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_653 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n7) );
  CMX2X1 U5 ( .A0(s4), .A1(s3), .S(n2), .Z(sum2[1]) );
  CMXI2X1 U6 ( .A0(n6), .A1(n4), .S(c_in2), .Z(n2) );
  CIVXL U7 ( .A(c_out01), .Z(n3) );
  CIVXL U8 ( .A(n3), .Z(n4) );
  CIVXL U9 ( .A(c_out00), .Z(n5) );
  CIVXL U10 ( .A(n5), .Z(n6) );
  CIVX1 U11 ( .A(c_out10), .Z(n9) );
  CIVX1 U12 ( .A(c_out11), .Z(n8) );
  CMXI2X1 U13 ( .A0(n8), .A1(n9), .S(n7), .Z(c_out2) );
  CMX2X1 U14 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module bit4_41 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_164 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_163 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_162 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_161 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(n7), .Z(n4) );
  CND2IX1 U4 ( .B(c_in4), .A(c_out400), .Z(n1) );
  CIVX1 U5 ( .A(s44[0]), .Z(n12) );
  CMXI2XL U6 ( .A0(n13), .A1(n12), .S(n7), .Z(sum4[2]) );
  CIVX1 U7 ( .A(s42[1]), .Z(n10) );
  CND2X1 U8 ( .A(c_out401), .B(c_in4), .Z(n2) );
  CND2X2 U9 ( .A(n1), .B(n2), .Z(n7) );
  CIVXL U10 ( .A(n4), .Z(n3) );
  CND2X2 U11 ( .A(n4), .B(c_out410), .Z(n5) );
  CND2X1 U12 ( .A(n7), .B(c_out411), .Z(n6) );
  CND2X2 U13 ( .A(n6), .B(n5), .Z(c_out4) );
  CMXI2XL U14 ( .A0(n15), .A1(n14), .S(n3), .Z(sum4[3]) );
  CIVX2 U15 ( .A(s41[0]), .Z(n9) );
  CIVX2 U16 ( .A(s42[0]), .Z(n8) );
  CMXI2X1 U17 ( .A0(n9), .A1(n8), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U18 ( .A(s41[1]), .Z(n11) );
  CMXI2X1 U19 ( .A0(n11), .A1(n10), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U20 ( .A(s43[0]), .Z(n13) );
  CIVX2 U21 ( .A(s43[1]), .Z(n15) );
  CIVX2 U22 ( .A(s44[1]), .Z(n14) );
endmodule


module Add_half_1313 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1314 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_657 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1314 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1313 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1315 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1316 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_658 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1316 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1315 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1317 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CNIVXL U2 ( .A(a), .Z(n2) );
  CEOXL U3 ( .A(b), .B(n2), .Z(sum) );
endmodule


module Add_half_1318 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_659 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1318 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1317 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1319 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1320 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_660 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1320 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1319 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_165 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_660 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_659 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_658 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_657 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2X1 U4 ( .A0(c_out11), .A1(c_out10), .S(n2), .Z(c_out2) );
  CMXI2XL U5 ( .A0(n6), .A1(n5), .S(n1), .Z(sum2[1]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX2 U7 ( .A(s1), .Z(n4) );
  CIVX2 U8 ( .A(s2), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module Add_half_1321 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1322 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_661 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1322 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1321 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1323 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1324 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_662 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1324 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1323 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1325 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n3;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
  CENXL U3 ( .A(n3), .B(a), .Z(sum) );
  CIVX2 U4 ( .A(b), .Z(n3) );
endmodule


module Add_half_1326 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_663 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1326 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1325 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1327 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1328 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_664 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1328 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1327 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_166 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_664 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_663 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_662 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_661 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2X1 U4 ( .A0(c_out11), .A1(c_out10), .S(n2), .Z(c_out2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module Add_half_1329 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1330 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_665 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1330 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1329 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1331 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1332 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_666 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1332 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1331 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1333 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CIVXL U3 ( .A(a), .Z(n2) );
  CIVX1 U4 ( .A(n2), .Z(n3) );
  CEOXL U5 ( .A(b), .B(n3), .Z(sum) );
endmodule


module Add_half_1334 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88962;
  assign c_out = net88962;

  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(net88962) );
endmodule


module Add_full_667 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1334 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1333 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1335 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CIVXL U3 ( .A(a), .Z(n2) );
  CIVXL U4 ( .A(n2), .Z(n3) );
  CEOXL U5 ( .A(b), .B(n3), .Z(sum) );
endmodule


module Add_half_1336 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88963, n1, n2, n3, n4;
  assign c_out = net88963;

  CND2X2 U1 ( .A(n3), .B(n4), .Z(sum) );
  CND2X2 U2 ( .A(n1), .B(b), .Z(n4) );
  CIVX2 U3 ( .A(a), .Z(n1) );
  CND2X1 U4 ( .A(a), .B(n2), .Z(n3) );
  CIVX1 U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(net88963) );
endmodule


module Add_full_668 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1336 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1335 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_167 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, net69579,
         net69580, net69578, n1, n2, n3, n4, n5;

  Add_full_668 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_667 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_666 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_665 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n2) );
  CNIVXL U4 ( .A(net69578), .Z(n1) );
  CIVX2 U5 ( .A(n3), .Z(net69578) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n3) );
  CMXI2X1 U7 ( .A0(net69579), .A1(net69580), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U8 ( .A0(n4), .A1(n5), .S(net69578), .Z(c_out2) );
  CIVX1 U9 ( .A(c_out11), .Z(n5) );
  CIVX2 U10 ( .A(c_out10), .Z(n4) );
  CIVX1 U11 ( .A(s2), .Z(net69580) );
  CIVX1 U12 ( .A(s1), .Z(net69579) );
  CMX2XL U13 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
endmodule


module Add_half_1337 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1338 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_669 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1338 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1337 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1339 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1340 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_670 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1340 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1339 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1341 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1342 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88964, n1, n2, n3, n4;
  assign c_out = net88964;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(net88964) );
endmodule


module Add_full_671 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1342 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1341 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1343 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CEOXL U2 ( .A(b), .B(n1), .Z(sum) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1344 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_672 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1344 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1343 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_168 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11;

  Add_full_672 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_671 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_670 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_669 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U4 ( .A(c_in2), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n3) );
  CIVX2 U6 ( .A(n3), .Z(n5) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n4) );
  CND2X2 U8 ( .A(c_out11), .B(n5), .Z(n6) );
  CND2X1 U9 ( .A(c_out10), .B(n4), .Z(n7) );
  CND2X2 U10 ( .A(n6), .B(n7), .Z(c_out2) );
  CMXI2X1 U11 ( .A0(n8), .A1(n9), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s1), .Z(n8) );
  CIVX2 U13 ( .A(s2), .Z(n9) );
  CMXI2XL U14 ( .A0(n11), .A1(n10), .S(n1), .Z(sum2[1]) );
  CIVX2 U15 ( .A(s3), .Z(n11) );
  CIVX2 U16 ( .A(s4), .Z(n10) );
endmodule


module bit4_42 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, net92553, net106504,
         net106503, net87626, net92984, n1, n2, n3, n4, n5, n6, n7;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_168 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_167 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_166 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_165 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(net92553), .Z(n5) );
  CND2X1 U4 ( .A(n6), .B(n7), .Z(sum4[2]) );
  CND2X1 U5 ( .A(c_out401), .B(c_in4), .Z(net92984) );
  CND2X2 U6 ( .A(net92984), .B(n2), .Z(net87626) );
  CIVX2 U7 ( .A(c_in4), .Z(n1) );
  CND2X2 U8 ( .A(c_out400), .B(n1), .Z(n2) );
  CND2XL U9 ( .A(c_out400), .B(n1), .Z(net106504) );
  CND2XL U10 ( .A(c_out401), .B(c_in4), .Z(net106503) );
  CMX2X1 U11 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U12 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMXI2X1 U13 ( .A0(n3), .A1(n4), .S(net87626), .Z(c_out4) );
  CIVX1 U14 ( .A(c_out411), .Z(n4) );
  CIVX1 U15 ( .A(c_out410), .Z(n3) );
  CND2X1 U16 ( .A(net106503), .B(net106504), .Z(net92553) );
  CND2X1 U17 ( .A(s44[0]), .B(net92553), .Z(n7) );
  CND2X1 U18 ( .A(s43[0]), .B(n5), .Z(n6) );
  CMX2X1 U19 ( .A0(s43[1]), .A1(s44[1]), .S(net92553), .Z(sum4[3]) );
endmodule


module Add_half_1345 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1346 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_673 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1346 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1345 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1347 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1348 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_674 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1348 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1347 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1349 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1350 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_675 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1350 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1349 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CND2X1 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_1351 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1352 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X2 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_676 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1352 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1351 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_169 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_676 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_675 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_674 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_673 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2XL U4 ( .A0(n7), .A1(n6), .S(n1), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n7) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
endmodule


module Add_half_1353 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
  CIVX2 U4 ( .A(b), .Z(n2) );
endmodule


module Add_half_1354 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_677 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1354 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1353 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1355 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1356 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_678 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1356 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1355 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1357 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1358 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_679 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1358 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1357 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_1359 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1360 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_680 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1360 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1359 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_170 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_680 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_679 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_678 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_677 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
endmodule


module Add_half_1361 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1362 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X2 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_681 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1362 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1361 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1363 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1364 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_682 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1364 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1363 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1365 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1366 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVX1 U1 ( .A(a), .Z(n1) );
  CND2X1 U2 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U3 ( .A(b), .Z(n2) );
  CND2XL U4 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U5 ( .A(n1), .B(b), .Z(n4) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_683 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1366 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1365 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1367 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1368 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_684 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1368 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1367 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_171 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_684 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_683 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_682 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_681 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMX2XL U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U5 ( .A(c_out10), .Z(n4) );
  CMXI2XL U6 ( .A0(n8), .A1(n7), .S(n1), .Z(sum2[1]) );
  CIVX2 U7 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX2 U9 ( .A(s1), .Z(n6) );
  CIVX2 U10 ( .A(s2), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s3), .Z(n8) );
  CIVX2 U13 ( .A(s4), .Z(n7) );
endmodule


module Add_half_1369 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1370 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_685 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1370 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1369 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1371 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1372 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_686 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1372 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1371 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1373 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1374 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_687 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1374 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1373 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1375 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1376 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_688 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1376 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1375 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_172 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_688 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_687 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_686 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_685 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CIVX20 U4 ( .A(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(c_out11), .Z(n3) );
  CIVX2 U6 ( .A(n2), .Z(n5) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(c_out10), .Z(n4) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(n5), .Z(c_out2) );
endmodule


module bit4_43 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_172 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_171 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_170 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_169 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(c_out411), .Z(n4) );
  CIVX2 U4 ( .A(c_in4), .Z(n1) );
  CMXI2X1 U5 ( .A0(c_out401), .A1(c_out400), .S(n1), .Z(n3) );
  CMX2XL U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CMX2X1 U7 ( .A0(s43[0]), .A1(s44[0]), .S(n2), .Z(sum4[2]) );
  CMXI2X1 U8 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out4) );
  CMX2XL U9 ( .A0(s43[1]), .A1(s44[1]), .S(n2), .Z(sum4[3]) );
  CMX2X1 U10 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U11 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX1 U12 ( .A(c_out410), .Z(n5) );
endmodule


module Add_half_1377 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1378 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_689 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1378 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1377 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1379 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1380 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CIVX2 U1 ( .A(b), .Z(n2) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_full_690 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1380 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1379 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1381 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1382 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n3), .B(n4), .Z(sum) );
  CND2X1 U3 ( .A(n1), .B(b), .Z(n4) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_691 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1382 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1381 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CND2X1 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_1383 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1384 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_692 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1384 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1383 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_173 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_692 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_691 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_690 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_689 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n2) );
  CMX2XL U4 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CMXI2X1 U5 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n3) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(c_out10), .Z(n5) );
  CIVX2 U10 ( .A(c_out11), .Z(n4) );
endmodule


module Add_half_1385 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1386 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_693 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1386 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1385 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1387 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_1388 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_694 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1388 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1387 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1389 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1390 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_695 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1390 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1389 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_1391 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1392 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_696 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1392 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1391 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_174 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_696 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_695 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_694 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_693 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_1393 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1394 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_697 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1394 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1393 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1395 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1396 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_698 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1396 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1395 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1397 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1398 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_699 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1398 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1397 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1399 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1400 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_700 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1400 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1399 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_175 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_700 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_699 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_698 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_697 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n5), .A1(n4), .S(n6), .Z(c_out2) );
  CIVX1 U4 ( .A(n3), .Z(n6) );
  CIVXL U5 ( .A(n6), .Z(n1) );
  CIVX1 U6 ( .A(n1), .Z(n2) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(c_out10), .Z(n5) );
  CIVX2 U10 ( .A(c_out11), .Z(n4) );
  CMXI2X1 U11 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
endmodule


module Add_half_1401 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1402 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_701 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1402 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1401 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1403 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1404 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_702 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1404 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1403 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1405 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1406 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_703 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1406 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1405 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1407 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1408 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_704 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1408 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1407 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_176 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_704 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_703 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_702 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_701 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CIVXL U4 ( .A(n6), .Z(n1) );
  CIVX1 U5 ( .A(n1), .Z(n2) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out10), .Z(n5) );
  CIVX2 U9 ( .A(c_out11), .Z(n4) );
  CIVX2 U10 ( .A(n3), .Z(n6) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(n6), .Z(c_out2) );
endmodule


module bit4_44 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_176 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_175 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_174 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_173 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVXL U4 ( .A(n1), .Z(n10) );
  CIVX1 U5 ( .A(s43[0]), .Z(n9) );
  CIVX1 U6 ( .A(c_out411), .Z(n2) );
  CIVX1 U7 ( .A(c_out410), .Z(n3) );
  CIVX1 U8 ( .A(s44[0]), .Z(n8) );
  CMXI2X1 U9 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out4) );
  CIVX2 U10 ( .A(s41[0]), .Z(n5) );
  CIVX2 U11 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U13 ( .A(s41[1]), .Z(n7) );
  CIVX2 U14 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U15 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CMXI2X1 U16 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CIVX2 U17 ( .A(s43[1]), .Z(n12) );
  CIVX2 U18 ( .A(s44[1]), .Z(n11) );
  CMXI2X1 U19 ( .A0(n12), .A1(n11), .S(n10), .Z(sum4[3]) );
endmodule


module bit8_11 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, net90172, net91740, net93721,
         net99223, net116545, net90171, n1, n2, n3, n4, n5, n6, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_44 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4({n11, b8[2:0]}), .c_in4(1'b0) );
  bit4_43 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4({n11, b8[2:0]}), .c_in4(1'b1) );
  bit4_42 A83 ( .sum4(s83), .c_out4(c_out810), .a4({a8[7], n8, n15, n16}), 
        .b4({b8[7:6], n10, b8[4]}), .c_in4(1'b0) );
  bit4_41 A84 ( .sum4(s84), .c_out4(c_out811), .a4({a8[7], n13, n15, n9}), 
        .b4({b8[7:6], n10, b8[4]}), .c_in4(1'b1) );
  CNIVX3 U3 ( .A(a8[4]), .Z(n9) );
  CIVX3 U4 ( .A(n1), .Z(sum8[2]) );
  CIVX2 U5 ( .A(n12), .Z(n13) );
  CMXI2X1 U6 ( .A0(s81[2]), .A1(s82[2]), .S(net90172), .Z(n1) );
  CIVX2 U7 ( .A(net90171), .Z(net90172) );
  CIVX3 U8 ( .A(n12), .Z(n8) );
  CMXI2X1 U9 ( .A0(n2), .A1(n3), .S(n4), .Z(c_out8) );
  CMXI2X1 U10 ( .A0(c_out801), .A1(c_out800), .S(net90171), .Z(n4) );
  CIVX2 U11 ( .A(c_in8), .Z(net90171) );
  CIVX1 U12 ( .A(c_out810), .Z(n3) );
  CIVX2 U13 ( .A(c_out811), .Z(n2) );
  CMXI2X1 U14 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(net93721) );
  CMXI2X1 U15 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(net116545) );
  CMX2X2 U16 ( .A0(s81[0]), .A1(s82[0]), .S(c_in8), .Z(sum8[0]) );
  CIVX1 U17 ( .A(a8[6]), .Z(n12) );
  CNIVX4 U18 ( .A(a8[4]), .Z(n16) );
  CIVX2 U19 ( .A(s83[2]), .Z(n17) );
  CND2X2 U20 ( .A(s84[0]), .B(net99223), .Z(n5) );
  CND2X1 U21 ( .A(s83[0]), .B(net93721), .Z(n6) );
  CND2X4 U22 ( .A(n5), .B(n6), .Z(sum8[4]) );
  CIVX1 U23 ( .A(net116545), .Z(net99223) );
  CMX2X2 U24 ( .A0(s84[1]), .A1(s83[1]), .S(net93721), .Z(sum8[5]) );
  CMX2X2 U25 ( .A0(s84[3]), .A1(s83[3]), .S(net91740), .Z(sum8[7]) );
  CMXI2X1 U26 ( .A0(n18), .A1(n17), .S(net116545), .Z(sum8[6]) );
  CNIVX1 U27 ( .A(net93721), .Z(net91740) );
  CIVX2 U28 ( .A(a8[5]), .Z(n14) );
  CNIVX4 U29 ( .A(b8[5]), .Z(n10) );
  CNIVX4 U30 ( .A(b8[3]), .Z(n11) );
  CMX2X1 U31 ( .A0(s81[3]), .A1(s82[3]), .S(net90172), .Z(sum8[3]) );
  CMX2X1 U32 ( .A0(s81[1]), .A1(s82[1]), .S(net90172), .Z(sum8[1]) );
  CIVX4 U33 ( .A(n14), .Z(n15) );
  CIVX1 U34 ( .A(s84[2]), .Z(n18) );
endmodule


module Add_half_1409 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1410 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_705 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1410 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1409 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1411 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1412 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_706 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1412 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1411 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1413 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1414 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_707 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1414 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1413 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1415 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1416 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_708 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1416 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1415 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_177 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_708 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_707 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_706 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_705 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2X1 U3 ( .A(c_out10), .B(n1), .Z(n2) );
  CND2X1 U4 ( .A(n2), .B(n3), .Z(c_out2) );
  CND2X1 U5 ( .A(c_out11), .B(n4), .Z(n3) );
  CIVX2 U6 ( .A(n4), .Z(n1) );
  CIVX1 U7 ( .A(n5), .Z(n4) );
  CIVXL U8 ( .A(n5), .Z(n8) );
  CMX2XL U9 ( .A0(s3), .A1(s4), .S(n8), .Z(sum2[1]) );
  CMXI2X1 U10 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n5) );
  CIVX2 U11 ( .A(s1), .Z(n7) );
  CIVX2 U12 ( .A(s2), .Z(n6) );
  CMXI2X1 U13 ( .A0(n7), .A1(n6), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_1417 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1418 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_709 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1418 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1417 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1419 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1420 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CNR2IXL U1 ( .B(a), .A(n2), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
  CIVXL U3 ( .A(b), .Z(n2) );
endmodule


module Add_full_710 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1420 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1419 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1421 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1422 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_711 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1422 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1421 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1423 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1424 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_712 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1424 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1423 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_178 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_712 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_711 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_710 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_709 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_1425 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1426 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_713 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1426 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1425 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1427 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CEOXL U2 ( .A(b), .B(n1), .Z(sum) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1428 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_714 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1428 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1427 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1429 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1430 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX1 U1 ( .A(n1), .B(a), .Z(sum) );
  CIVXL U2 ( .A(b), .Z(n1) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_715 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1430 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1429 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1431 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1432 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX1 U1 ( .A(n1), .B(a), .Z(sum) );
  CIVXL U2 ( .A(b), .Z(n1) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_716 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1432 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1431 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_179 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_716 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_715 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_714 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_713 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s2), .Z(n4) );
  CIVX1 U4 ( .A(s1), .Z(n5) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n6) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_1433 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1434 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_717 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1434 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1433 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1435 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOX1 U1 ( .A(b), .B(n1), .Z(sum) );
  CNIVXL U2 ( .A(a), .Z(n1) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1436 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_718 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1436 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1435 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1437 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1438 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_719 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1438 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1437 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1439 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1440 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_720 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1440 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1439 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_180 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_720 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_719 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_718 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_717 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2XL U4 ( .A0(n7), .A1(n6), .S(n5), .Z(sum2[1]) );
  CIVX1 U5 ( .A(n2), .Z(n5) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CIVX1 U7 ( .A(s4), .Z(n6) );
  CIVX1 U8 ( .A(s3), .Z(n7) );
  CMX2X1 U9 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U10 ( .A(c_out10), .Z(n4) );
  CIVX2 U11 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U12 ( .A0(n4), .A1(n3), .S(n5), .Z(c_out2) );
endmodule


module bit4_45 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_180 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_179 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_178 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_177 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2XL U4 ( .A0(n6), .A1(n5), .S(n4), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMXI2X1 U6 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out4) );
  CIVX1 U7 ( .A(n1), .Z(n4) );
  CMX2X1 U8 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U9 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX1 U10 ( .A(c_out410), .Z(n3) );
  CIVX2 U11 ( .A(c_out411), .Z(n2) );
  CIVX2 U12 ( .A(s43[1]), .Z(n6) );
  CIVX2 U13 ( .A(s44[1]), .Z(n5) );
endmodule


module Add_half_1441 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1442 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_721 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1442 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1441 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1443 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1444 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX2 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_722 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1444 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1443 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1445 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1446 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_723 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1446 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1445 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1447 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1448 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_724 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1448 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1447 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_181 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_724 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_723 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_722 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_721 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s3), .Z(n4) );
  CIVX2 U9 ( .A(s4), .Z(n3) );
endmodule


module Add_half_1449 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1450 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_725 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1450 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1449 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1451 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1452 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_726 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1452 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1451 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1453 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1454 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_727 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1454 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1453 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1455 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1456 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_728 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1456 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1455 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_182 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_728 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_727 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_726 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_725 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_1457 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1458 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_729 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1458 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1457 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1459 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1460 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_730 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1460 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1459 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1461 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1462 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_731 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1462 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1461 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1463 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1464 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX1 U1 ( .A(a), .B(n1), .Z(sum) );
  CIVXL U2 ( .A(b), .Z(n1) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_732 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1464 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1463 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_183 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_732 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_731 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_730 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_729 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n4) );
endmodule


module Add_half_1465 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1466 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_733 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1466 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1465 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1467 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1468 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_734 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1468 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1467 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1469 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1470 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX1 U1 ( .A(a), .B(n1), .Z(sum) );
  CIVXL U2 ( .A(b), .Z(n1) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_735 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1470 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1469 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1471 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1472 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX1 U1 ( .A(a), .B(n1), .Z(sum) );
  CIVXL U2 ( .A(b), .Z(n1) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_736 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1472 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1471 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_184 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_736 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_735 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_734 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_733 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_46 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_184 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_183 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_182 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_181 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(n10), .A1(n9), .S(n11), .Z(sum4[2]) );
  CMXI2XL U4 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U5 ( .A(c_out411), .Z(n3) );
  CMXI2X1 U6 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out4) );
  CIVX1 U7 ( .A(n1), .Z(n11) );
  CIVX2 U8 ( .A(c_out410), .Z(n4) );
  CIVX1 U9 ( .A(s42[0]), .Z(n5) );
  CIVX1 U10 ( .A(s41[0]), .Z(n6) );
  CMX2XL U11 ( .A0(s43[1]), .A1(s44[1]), .S(n11), .Z(sum4[3]) );
  CMXI2X1 U12 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CMXI2X1 U13 ( .A0(n6), .A1(n5), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U14 ( .A(s41[1]), .Z(n8) );
  CIVX2 U15 ( .A(s42[1]), .Z(n7) );
  CMXI2X1 U16 ( .A0(n8), .A1(n7), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U17 ( .A(s43[0]), .Z(n10) );
  CIVX2 U18 ( .A(s44[0]), .Z(n9) );
endmodule


module Add_half_1473 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1474 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_737 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1474 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1473 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1475 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1476 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_738 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1476 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1475 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1477 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1478 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_739 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1478 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1477 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1479 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1480 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_740 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1480 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1479 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_185 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_740 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_739 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_738 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_737 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_1481 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1482 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_741 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1482 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1481 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1483 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1484 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_742 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1484 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1483 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1485 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1486 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_743 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1486 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1485 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1487 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1488 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_744 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1488 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1487 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_186 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_744 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_743 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_742 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_741 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CIVX2 U7 ( .A(s1), .Z(n3) );
  CIVX2 U8 ( .A(s2), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_1489 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1490 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_745 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1490 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1489 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1491 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1492 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_746 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1492 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1491 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1493 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1494 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_747 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1494 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1493 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1495 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1496 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_748 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1496 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1495 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_187 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_748 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_747 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_746 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_745 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module Add_half_1497 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1498 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_749 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1498 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1497 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1499 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1500 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_750 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1500 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1499 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1501 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1502 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_751 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1502 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1501 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1503 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1504 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_752 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1504 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1503 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_188 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_752 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_751 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_750 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_749 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module bit4_47 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_188 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_187 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_186 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_185 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n7), .Z(sum4[0]) );
  CMX2XL U3 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U4 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U5 ( .A(c_out410), .Z(n3) );
  CIVX2 U6 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
  CIVX2 U11 ( .A(s43[1]), .Z(n6) );
  CIVX2 U12 ( .A(s44[1]), .Z(n5) );
  CMXI2X1 U13 ( .A0(n6), .A1(n5), .S(n4), .Z(sum4[3]) );
  CIVX2 U14 ( .A(c_in4), .Z(n7) );
endmodule


module Add_half_1505 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1506 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_753 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1506 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1505 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1507 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1508 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_754 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1508 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1507 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1509 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1510 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_755 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1510 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1509 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1511 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1512 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_756 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1512 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1511 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_189 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_756 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_755 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_754 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_753 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U7 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_1513 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1514 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_757 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1514 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1513 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1515 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1516 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_758 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1516 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1515 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1517 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1518 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_759 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1518 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1517 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1519 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1520 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_760 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1520 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1519 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_190 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_760 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_759 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_758 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_757 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_1521 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1522 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_761 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1522 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1521 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1523 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1524 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_762 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1524 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1523 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1525 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1526 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_763 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1526 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1525 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1527 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1528 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_764 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1528 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1527 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_191 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_764 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_763 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_762 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_761 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_1529 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1530 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_765 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1530 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1529 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1531 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1532 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_766 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1532 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1531 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1533 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1534 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_767 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1534 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1533 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1535 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1536 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_768 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1536 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1535 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_192 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_768 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_767 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_766 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_765 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module bit4_48 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_192 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_191 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_190 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_189 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n9), .Z(sum4[0]) );
  CIVX2 U3 ( .A(c_out410), .Z(n3) );
  CMX2XL U4 ( .A0(s43[1]), .A1(s44[1]), .S(n8), .Z(sum4[3]) );
  CIVX1 U5 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n8) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U10 ( .A(s41[1]), .Z(n5) );
  CIVX2 U11 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U13 ( .A(s43[0]), .Z(n7) );
  CIVX2 U14 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U15 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX2 U16 ( .A(c_in4), .Z(n9) );
endmodule


module bit8_12 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   n14, c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n6, n7,
         n8, n9, n10, n11, n12, n13;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_48 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_47 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_46 A83 ( .sum4(s83), .c_out4(c_out810), .a4({a8[7], n10, a8[5], n7}), 
        .b4(b8[7:4]), .c_in4(1'b0) );
  bit4_45 A84 ( .sum4(s84), .c_out4(c_out811), .a4({a8[7], n10, a8[5], n9}), 
        .b4(b8[7:4]), .c_in4(1'b1) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n13), .Z(sum8[0]) );
  CND2X1 U3 ( .A(c_out810), .B(n1), .Z(n2) );
  CND2X1 U4 ( .A(c_out811), .B(n12), .Z(n3) );
  CND2X2 U5 ( .A(n2), .B(n3), .Z(c_out8) );
  CIVX1 U6 ( .A(n12), .Z(n1) );
  CMX2X2 U7 ( .A0(s83[3]), .A1(s84[3]), .S(n6), .Z(sum8[7]) );
  CIVX3 U8 ( .A(n14), .Z(n4) );
  CIVX4 U9 ( .A(n4), .Z(sum8[6]) );
  CMX2X1 U10 ( .A0(s83[2]), .A1(s84[2]), .S(n6), .Z(n14) );
  CMX2X2 U11 ( .A0(s83[1]), .A1(s84[1]), .S(n6), .Z(sum8[5]) );
  CMX2X2 U12 ( .A0(s83[0]), .A1(s84[0]), .S(n12), .Z(sum8[4]) );
  CIVX2 U14 ( .A(n11), .Z(n12) );
  CNIVX4 U15 ( .A(n12), .Z(n6) );
  CIVX3 U16 ( .A(n8), .Z(n7) );
  CIVX3 U17 ( .A(n8), .Z(n9) );
  CIVX2 U18 ( .A(a8[4]), .Z(n8) );
  CNIVX4 U19 ( .A(a8[6]), .Z(n10) );
  CMX2X2 U20 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2X2 U21 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2X2 U22 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMXI2X1 U23 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n11) );
  CIVX2 U24 ( .A(c_in8), .Z(n13) );
endmodule


module bit32_3 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   c1, c2, c3, n1, n2, n3, n4, n5;

  bit8_12 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8(a32[7:0]), .b8(b32[7:0]), 
        .c_in8(c_in32) );
  bit8_11 A322 ( .sum8(sum32[15:8]), .c_out8(c2), .a8({a32[15:9], n3}), .b8(
        b32[15:8]), .c_in8(c1) );
  bit8_10 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8({a32[23], n1, 
        a32[21:17], n5}), .b8(b32[23:16]), .c_in8(c2) );
  bit8_9 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8(a32[31:24]), .b8(
        b32[31:24]), .c_in8(c3) );
  CNIVX4 U1 ( .A(a32[22]), .Z(n1) );
  CIVX2 U2 ( .A(a32[8]), .Z(n2) );
  CIVX4 U3 ( .A(n2), .Z(n3) );
  CIVX2 U4 ( .A(a32[16]), .Z(n4) );
  CIVX4 U5 ( .A(n4), .Z(n5) );
endmodule


module Add_half_1537 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1538 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_769 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1538 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1537 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1539 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1540 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_770 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1540 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1539 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1541 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1542 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_771 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1542 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1541 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1543 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1544 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_772 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1544 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1543 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_193 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_772 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_771 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_770 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_769 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1545 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1546 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_773 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1546 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1545 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1547 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1548 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_774 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1548 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1547 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1549 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1550 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_775 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1550 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1549 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1551 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1552 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_776 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1552 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1551 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_194 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_776 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_775 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_774 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_773 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1553 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1554 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_777 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1554 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1553 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1555 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1556 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_778 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1556 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1555 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1557 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1558 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_779 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1558 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1557 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1559 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1560 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_780 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1560 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1559 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_195 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_780 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_779 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_778 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_777 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_1561 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1562 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_781 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1562 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1561 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1563 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1564 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_782 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1564 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1563 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1565 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1566 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_783 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1566 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1565 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1567 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1568 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_784 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1568 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1567 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_196 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_784 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_783 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_782 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_781 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s3), .Z(n6) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module bit4_49 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_196 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_195 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_194 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_193 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U6 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2X1 U7 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
endmodule


module Add_half_1569 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1570 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_785 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1570 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1569 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1571 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1572 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_786 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1572 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1571 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1573 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1574 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_787 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1574 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1573 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1575 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1576 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_788 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1576 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1575 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_197 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_788 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_787 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_786 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_785 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1577 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1578 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_789 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1578 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1577 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1579 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1580 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_790 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1580 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1579 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1581 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1582 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_791 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1582 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1581 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1583 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1584 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_792 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1584 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1583 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_198 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_792 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_791 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_790 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_789 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1585 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1586 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_793 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1586 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1585 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1587 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1588 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_794 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1588 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1587 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1589 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1590 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_795 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1590 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1589 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1591 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1592 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_796 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1592 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1591 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_199 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_796 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_795 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_794 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_793 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_1593 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1594 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_797 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1594 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1593 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1595 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1596 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_798 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1596 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1595 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1597 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1598 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_799 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1598 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1597 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1599 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1600 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_800 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1600 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1599 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_200 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_800 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_799 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_798 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_797 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n4) );
endmodule


module bit4_50 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_200 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_199 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_198 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_197 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n9), .A1(n8), .S(n1), .Z(sum4[3]) );
  CMX2X2 U4 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMX2X1 U5 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CIVX2 U6 ( .A(s41[0]), .Z(n3) );
  CIVX2 U7 ( .A(s42[0]), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U9 ( .A(s41[1]), .Z(n5) );
  CIVX2 U10 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(s43[0]), .Z(n7) );
  CIVX2 U13 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n1), .Z(sum4[2]) );
  CIVX2 U15 ( .A(s43[1]), .Z(n9) );
  CIVX2 U16 ( .A(s44[1]), .Z(n8) );
endmodule


module Add_half_1601 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1602 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_801 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1602 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1601 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1603 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1604 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_802 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1604 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1603 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1605 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1606 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_803 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1606 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1605 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1607 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1608 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_804 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1608 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1607 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_201 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_804 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_803 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_802 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_801 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(n1), .Z(n4) );
  CIVX2 U6 ( .A(s1), .Z(n3) );
  CIVX2 U7 ( .A(s2), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_1609 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1610 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_805 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1610 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1609 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1611 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1612 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_806 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1612 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1611 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1613 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1614 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_807 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1614 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1613 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1615 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1616 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_808 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1616 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1615 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_202 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_808 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_807 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_806 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_805 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U7 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_1617 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1618 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_809 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1618 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1617 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1619 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1620 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_810 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1620 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1619 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1621 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1622 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_811 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1622 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1621 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1623 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1624 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_812 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1624 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1623 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_203 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_812 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_811 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_810 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_809 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_1625 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1626 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_813 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1626 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1625 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1627 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1628 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_814 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1628 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1627 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1629 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1630 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_815 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1630 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1629 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1631 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1632 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_816 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1632 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1631 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_204 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_816 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_815 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_814 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_813 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_51 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_204 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_203 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_202 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_201 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U4 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n4) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
  CIVX2 U11 ( .A(s43[1]), .Z(n6) );
  CIVX2 U12 ( .A(s44[1]), .Z(n5) );
  CMXI2X1 U13 ( .A0(n6), .A1(n5), .S(n4), .Z(sum4[3]) );
endmodule


module Add_half_1633 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1634 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_817 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1634 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1633 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1635 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1636 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_818 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1636 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1635 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1637 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1638 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_819 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1638 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1637 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1639 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1640 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_820 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1640 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1639 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_205 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_820 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_819 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_818 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_817 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(s3), .Z(n3) );
  CIVX2 U8 ( .A(s4), .Z(n2) );
endmodule


module Add_half_1641 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1642 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_821 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1642 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1641 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1643 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1644 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_822 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1644 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1643 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1645 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1646 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_823 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1646 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1645 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1647 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1648 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_824 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1648 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1647 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_206 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_824 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_823 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_822 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_821 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s3), .Z(n4) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_1649 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1650 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_825 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1650 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1649 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1651 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1652 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_826 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1652 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1651 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1653 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1654 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_827 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1654 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1653 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1655 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1656 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_828 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1656 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1655 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_207 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_828 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_827 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_826 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_825 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_1657 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1658 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_829 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1658 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1657 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1659 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1660 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_830 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1660 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1659 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1661 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1662 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_831 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1662 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1661 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1663 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1664 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_832 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1664 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1663 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_208 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_832 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_831 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_830 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_829 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module bit4_52 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_208 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_207 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_206 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_205 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out4) );
  CMX2XL U4 ( .A0(s43[1]), .A1(s44[1]), .S(n6), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n6) );
  CIVX2 U11 ( .A(s43[0]), .Z(n5) );
  CIVX2 U12 ( .A(s44[0]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(n6), .Z(sum4[2]) );
endmodule


module bit8_13 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_52 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_51 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_50 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_49 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2XL U3 ( .A0(s83[3]), .A1(s84[3]), .S(n1), .Z(sum8[7]) );
  CMXI2XL U4 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out8) );
  CMX2X2 U5 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMXI2XL U6 ( .A0(n7), .A1(n6), .S(c_in8), .Z(sum8[1]) );
  CMX2X1 U7 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CIVX2 U8 ( .A(s81[1]), .Z(n7) );
  CMX2X2 U9 ( .A0(s83[0]), .A1(s84[0]), .S(n1), .Z(sum8[4]) );
  CMX2X1 U10 ( .A0(s83[2]), .A1(s84[2]), .S(n1), .Z(sum8[6]) );
  CIVX1 U11 ( .A(s82[0]), .Z(n4) );
  CMX2X1 U12 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2X1 U13 ( .A0(s83[1]), .A1(s84[1]), .S(n1), .Z(sum8[5]) );
  CIVX2 U14 ( .A(c_out810), .Z(n3) );
  CIVX2 U15 ( .A(c_out811), .Z(n2) );
  CIVX2 U16 ( .A(s81[0]), .Z(n5) );
  CMXI2X1 U17 ( .A0(n5), .A1(n4), .S(c_in8), .Z(sum8[0]) );
  CIVX2 U18 ( .A(s82[1]), .Z(n6) );
endmodule


module Add_half_1665 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1666 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_833 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1666 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1665 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1667 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1668 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_834 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1668 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1667 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1669 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1670 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_835 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1670 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1669 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1671 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1672 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_836 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1672 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1671 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_209 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_836 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_835 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_834 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_833 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n7), .A1(n6), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n7) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
endmodule


module Add_half_1673 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1674 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_837 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1674 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1673 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1675 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1676 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_838 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1676 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1675 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1677 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1678 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_839 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1678 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1677 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1679 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1680 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_840 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1680 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1679 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_210 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_840 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_839 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_838 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_837 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(s3), .Z(n4) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_1681 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1682 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_841 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1682 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1681 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1683 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1684 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_842 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1684 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1683 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1685 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1686 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_843 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1686 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1685 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1687 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1688 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_844 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1688 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1687 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_211 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_844 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_843 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_842 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_841 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(n1), .Z(n6) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s3), .Z(n8) );
  CIVX2 U13 ( .A(s4), .Z(n7) );
endmodule


module Add_half_1689 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1690 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_845 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1690 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1689 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1691 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1692 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_846 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1692 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1691 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1693 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1694 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_847 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1694 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1693 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1695 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1696 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_848 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1696 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1695 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_212 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_848 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_847 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_846 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_845 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2XL U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX1 U5 ( .A(n1), .Z(n4) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_53 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_212 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_211 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_210 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_209 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n2), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n2), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(c_out410), .A1(c_out411), .S(n2), .Z(c_out4) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U7 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n2) );
endmodule


module Add_half_1697 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1698 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_849 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1698 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1697 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1699 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1700 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_850 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1700 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1699 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1701 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1702 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_851 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1702 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1701 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1703 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1704 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_852 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1704 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1703 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_213 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_852 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_851 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_850 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_849 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_1705 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1706 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_853 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1706 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1705 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1707 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1708 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_854 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1708 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1707 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1709 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1710 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_855 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1710 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1709 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1711 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1712 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_856 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1712 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1711 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_214 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_856 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_855 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_854 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_853 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_1713 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1714 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_857 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1714 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1713 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1715 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1716 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_858 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1716 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1715 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1717 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1718 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_859 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1718 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1717 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1719 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1720 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_860 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1720 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1719 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_215 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_860 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_859 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_858 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_857 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_1721 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1722 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_861 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1722 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1721 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1723 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1724 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_862 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1724 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1723 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1725 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1726 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_863 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1726 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1725 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1727 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1728 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_864 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1728 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1727 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_216 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_864 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_863 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_862 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_861 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_54 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_216 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_215 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_214 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_213 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n11), .A1(n10), .S(n1), .Z(sum4[3]) );
  CMXI2XL U4 ( .A0(n9), .A1(n8), .S(n1), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out4) );
  CIVX2 U9 ( .A(s41[0]), .Z(n5) );
  CIVX2 U10 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U12 ( .A(s41[1]), .Z(n7) );
  CIVX2 U13 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U15 ( .A(s43[0]), .Z(n9) );
  CIVX2 U16 ( .A(s44[0]), .Z(n8) );
  CIVX2 U17 ( .A(s43[1]), .Z(n11) );
  CIVX2 U18 ( .A(s44[1]), .Z(n10) );
endmodule


module Add_half_1729 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1730 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_865 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1730 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1729 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1731 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1732 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_866 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1732 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1731 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1733 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1734 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_867 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1734 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1733 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1735 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1736 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_868 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1736 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1735 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_217 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_868 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_867 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_866 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_865 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_1737 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1738 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_869 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1738 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1737 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1739 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1740 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_870 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1740 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1739 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1741 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1742 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_871 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1742 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1741 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1743 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1744 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_872 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1744 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1743 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_218 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_872 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_871 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_870 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_869 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(s3), .Z(n6) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_1745 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1746 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_873 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1746 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1745 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1747 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1748 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_874 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1748 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1747 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1749 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1750 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_875 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1750 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1749 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1751 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1752 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_876 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1752 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1751 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_219 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_876 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_875 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_874 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_873 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_1753 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_1754 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_877 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1754 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1753 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1755 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1756 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_878 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1756 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1755 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1757 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1758 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_879 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_1758 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1757 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1759 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1760 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_880 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1760 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1759 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_220 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_880 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_879 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_878 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_877 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_55 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_220 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_219 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_218 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_217 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n8), .Z(sum4[3]) );
  CMX2X1 U4 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U5 ( .A(c_out410), .Z(n3) );
  CIVX2 U6 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n8) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U10 ( .A(s41[0]), .Z(n5) );
  CIVX2 U11 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U13 ( .A(s43[0]), .Z(n7) );
  CIVX2 U14 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U15 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
endmodule


module Add_half_1761 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1762 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_881 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1762 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1761 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1763 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1764 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_882 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1764 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1763 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1765 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1766 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_883 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1766 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1765 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1767 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1768 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_884 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1768 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1767 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_221 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_884 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_883 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_882 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_881 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_1769 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1770 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_885 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1770 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1769 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1771 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1772 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_886 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1772 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1771 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1773 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1774 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_887 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1774 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1773 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1775 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1776 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_888 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1776 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1775 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_222 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_888 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_887 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_886 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_885 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_1777 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1778 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_889 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1778 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1777 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1779 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1780 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_890 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1780 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1779 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1781 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1782 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_891 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1782 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1781 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1783 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1784 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_892 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1784 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1783 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_223 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_892 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_891 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_890 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_889 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_1785 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1786 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_893 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1786 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1785 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1787 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1788 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_894 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1788 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1787 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1789 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(a), .B(n2), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_1790 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_895 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1790 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1789 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1791 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1792 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_896 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1792 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1791 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_224 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_896 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_895 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_894 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_893 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_56 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_224 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_223 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_222 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_221 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(c_in4), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out401), .A1(c_out400), .S(n1), .Z(n2) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U6 ( .A(c_out410), .Z(n4) );
  CIVX2 U7 ( .A(c_out411), .Z(n3) );
  CIVX2 U8 ( .A(n2), .Z(n9) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n9), .Z(c_out4) );
  CIVX2 U10 ( .A(s41[1]), .Z(n6) );
  CIVX2 U11 ( .A(s42[1]), .Z(n5) );
  CMXI2X1 U12 ( .A0(n6), .A1(n5), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U13 ( .A(s43[0]), .Z(n8) );
  CIVX2 U14 ( .A(s44[0]), .Z(n7) );
  CMXI2X1 U15 ( .A0(n8), .A1(n7), .S(n9), .Z(sum4[2]) );
  CIVX2 U16 ( .A(s43[1]), .Z(n11) );
  CIVX2 U17 ( .A(s44[1]), .Z(n10) );
  CMXI2X1 U18 ( .A0(n11), .A1(n10), .S(n9), .Z(sum4[3]) );
endmodule


module bit8_14 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_56 A81 ( .sum4(s81), .c_out4(c_out800), .a4({a8[3:1], n6}), .b4({n5, 
        b8[2:1], n2}), .c_in4(1'b0) );
  bit4_55 A82 ( .sum4(s82), .c_out4(c_out801), .a4({a8[3:1], n4}), .b4({n5, 
        b8[2:1], n2}), .c_in4(1'b1) );
  bit4_54 A83 ( .sum4(s83), .c_out4(c_out810), .a4({a8[7:5], n3}), .b4(b8[7:4]), .c_in4(1'b0) );
  bit4_53 A84 ( .sum4(s84), .c_out4(c_out811), .a4({a8[7:5], n3}), .b4(b8[7:4]), .c_in4(1'b1) );
  CNIVX1 U3 ( .A(c_in8), .Z(n1) );
  CMX2X1 U4 ( .A0(c_out810), .A1(c_out811), .S(n12), .Z(c_out8) );
  CIVX2 U5 ( .A(n7), .Z(n12) );
  CNIVX4 U6 ( .A(b8[0]), .Z(n2) );
  CMX2X2 U7 ( .A0(s83[2]), .A1(s84[2]), .S(n12), .Z(sum8[6]) );
  CNIVX4 U8 ( .A(a8[4]), .Z(n3) );
  CMXI2X4 U9 ( .A0(n11), .A1(n10), .S(n12), .Z(sum8[4]) );
  CNIVX4 U10 ( .A(a8[0]), .Z(n4) );
  CNIVX4 U11 ( .A(b8[3]), .Z(n5) );
  CNIVX4 U12 ( .A(a8[0]), .Z(n6) );
  CMX2X1 U13 ( .A0(s81[3]), .A1(s82[3]), .S(n1), .Z(sum8[3]) );
  CMX2X1 U14 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2X1 U15 ( .A0(s83[3]), .A1(s84[3]), .S(n12), .Z(sum8[7]) );
  CMX2X1 U16 ( .A0(s83[1]), .A1(s84[1]), .S(n12), .Z(sum8[5]) );
  CMXI2X2 U17 ( .A0(n9), .A1(n8), .S(c_in8), .Z(sum8[0]) );
  CMX2X1 U18 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMXI2X1 U19 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n7) );
  CIVX2 U20 ( .A(s81[0]), .Z(n9) );
  CIVX2 U21 ( .A(s82[0]), .Z(n8) );
  CIVX2 U22 ( .A(s83[0]), .Z(n11) );
  CIVX2 U23 ( .A(s84[0]), .Z(n10) );
endmodule


module Add_half_1793 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1794 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_897 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1794 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1793 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1795 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1796 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_898 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1796 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1795 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1797 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1798 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_899 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1798 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1797 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1799 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1800 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_900 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1800 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1799 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_225 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_900 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_899 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_898 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_897 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_1801 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1802 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_901 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1802 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1801 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1803 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1804 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_902 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1804 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1803 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1805 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1806 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_903 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1806 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1805 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1807 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1808 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_904 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1808 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1807 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_226 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_904 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_903 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_902 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_901 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_1809 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1810 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_905 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1810 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1809 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1811 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1812 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_906 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1812 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1811 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1813 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1814 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_907 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1814 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1813 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1815 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1816 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_908 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1816 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1815 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_227 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_908 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_907 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_906 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_905 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U4 ( .A(s3), .Z(n5) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(s4), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module Add_half_1817 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1818 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_909 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1818 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1817 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1819 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1820 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_910 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1820 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1819 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1821 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1822 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_911 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1822 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1821 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1823 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1824 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_912 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1824 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1823 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_228 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_912 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_911 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_910 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_909 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVXL U4 ( .A(s3), .Z(n5) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(s4), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module bit4_57 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_228 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_227 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_226 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_225 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n7), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n7), .Z(sum4[0]) );
  CMX2X1 U3 ( .A0(c_out410), .A1(c_out411), .S(n4), .Z(c_out4) );
  CMXI2X1 U4 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U5 ( .A(n1), .Z(n4) );
  CIVX2 U6 ( .A(s43[0]), .Z(n3) );
  CIVX2 U7 ( .A(s44[0]), .Z(n2) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n4), .Z(sum4[2]) );
  CIVX2 U11 ( .A(s43[1]), .Z(n6) );
  CIVX2 U12 ( .A(s44[1]), .Z(n5) );
  CMXI2X1 U13 ( .A0(n6), .A1(n5), .S(n4), .Z(sum4[3]) );
  CIVX2 U14 ( .A(c_in4), .Z(n7) );
endmodule


module Add_half_1825 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1826 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_913 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1826 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1825 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1827 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1828 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_914 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1828 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1827 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1829 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1830 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_915 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1830 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1829 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1831 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1832 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_916 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1832 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1831 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_229 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_916 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_915 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_914 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_913 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U7 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_1833 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1834 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_917 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1834 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1833 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1835 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1836 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_918 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1836 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1835 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1837 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1838 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_919 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1838 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1837 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_1839 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_1840 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_920 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_1840 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1839 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_230 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_920 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_919 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_918 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_917 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s3), .Z(n4) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_1841 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1842 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_921 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1842 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1841 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1843 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1844 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_922 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1844 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1843 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1845 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1846 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_923 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1846 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1845 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1847 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1848 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_924 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1848 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1847 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_231 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_924 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_923 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_922 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_921 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVXL U5 ( .A(s3), .Z(n5) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module Add_half_1849 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1850 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_925 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1850 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1849 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1851 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1852 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_926 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1852 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1851 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1853 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_1854 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_927 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1854 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1853 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_1855 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1856 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_928 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1856 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1855 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_232 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_928 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_927 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_926 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_925 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U8 ( .A(s3), .Z(n5) );
  CIVX2 U9 ( .A(s4), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module bit4_58 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_232 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_231 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_230 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_229 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n7), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n7), .Z(sum4[0]) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n6), .Z(sum4[3]) );
  CIVX1 U4 ( .A(c_out411), .Z(n2) );
  CIVX1 U5 ( .A(c_out410), .Z(n3) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out4) );
  CIVX2 U11 ( .A(s43[0]), .Z(n5) );
  CIVX2 U12 ( .A(s44[0]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(n6), .Z(sum4[2]) );
  CIVX2 U14 ( .A(c_in4), .Z(n7) );
endmodule


module Add_half_1857 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1858 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_929 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1858 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1857 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1859 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1860 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_930 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1860 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1859 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1861 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1862 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_931 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1862 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1861 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1863 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1864 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_932 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1864 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1863 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_233 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_932 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_931 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_930 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_929 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1865 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1866 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_933 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1866 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1865 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1867 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1868 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_934 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1868 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1867 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1869 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1870 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_935 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1870 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1869 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1871 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1872 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_936 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1872 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1871 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_234 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_936 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_935 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_934 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_933 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1873 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1874 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_937 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1874 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1873 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1875 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1876 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_938 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1876 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1875 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1877 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1878 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_939 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1878 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1877 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1879 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1880 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_940 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1880 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1879 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_235 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_940 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_939 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_938 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_937 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1881 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1882 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_941 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1882 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1881 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1883 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1884 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_942 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1884 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1883 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1885 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1886 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_943 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1886 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1885 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1887 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1888 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_944 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1888 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1887 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_236 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_944 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_943 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_942 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_941 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_59 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_236 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_235 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_234 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_233 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_1889 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1890 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_945 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1890 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1889 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1891 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1892 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_946 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1892 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1891 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1893 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1894 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_947 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1894 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1893 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1895 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1896 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_948 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1896 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1895 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_237 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_948 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_947 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_946 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_945 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1897 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1898 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_949 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1898 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1897 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1899 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1900 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_950 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1900 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1899 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1901 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1902 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_951 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1902 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1901 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1903 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1904 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_952 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1904 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1903 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_238 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_952 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_951 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_950 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_949 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1905 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1906 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_953 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1906 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1905 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1907 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1908 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_954 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1908 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1907 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1909 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1910 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_955 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1910 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1909 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1911 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1912 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_956 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1912 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1911 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_239 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_956 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_955 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_954 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_953 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1913 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1914 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_957 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1914 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1913 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1915 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1916 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_958 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1916 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1915 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1917 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1918 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_959 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1918 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1917 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1919 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1920 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_960 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1920 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1919 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_240 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_960 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_959 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_958 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_957 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_60 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_240 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_239 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_238 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_237 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_15 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n2, n3, n4;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_60 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_59 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_58 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_57 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n4), .C(s83[1]), .D(n2), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n4), .C(s83[0]), .D(n2), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n3), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n3), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n3), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n3), .Z(sum8[0]) );
  CMX2X2 U3 ( .A0(s84[2]), .A1(s83[2]), .S(n2), .Z(sum8[6]) );
  CMX2X1 U4 ( .A0(c_out810), .A1(c_out811), .S(n4), .Z(c_out8) );
  CMX2X2 U5 ( .A0(s83[3]), .A1(s84[3]), .S(n4), .Z(sum8[7]) );
  CMXI2X1 U6 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n2) );
  CIVX2 U7 ( .A(n2), .Z(n4) );
  CIVX2 U14 ( .A(c_in8), .Z(n3) );
endmodule


module Add_half_1921 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1922 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_961 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1922 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1921 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1923 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1924 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_962 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1924 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1923 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1925 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1926 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_963 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1926 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1925 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1927 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1928 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_964 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1928 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1927 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_241 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_964 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_963 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_962 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_961 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1929 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1930 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_965 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1930 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1929 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1931 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1932 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_966 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1932 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1931 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1933 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1934 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_967 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1934 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1933 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1935 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1936 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_968 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1936 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1935 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_242 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_968 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_967 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_966 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_965 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1937 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1938 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_969 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1938 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1937 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1939 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1940 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_970 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1940 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1939 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1941 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1942 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_971 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1942 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1941 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1943 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1944 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_972 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1944 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1943 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_243 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_972 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_971 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_970 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_969 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1945 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1946 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_973 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1946 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1945 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1947 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1948 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_974 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1948 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1947 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1949 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1950 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_975 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1950 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1949 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1951 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1952 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_976 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1952 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1951 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_244 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_976 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_975 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_974 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_973 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_61 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_244 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_243 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_242 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_241 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_1953 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1954 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_977 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1954 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1953 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1955 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1956 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_978 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1956 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1955 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1957 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1958 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_979 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1958 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1957 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1959 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1960 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_980 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1960 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1959 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_245 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_980 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_979 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_978 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_977 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1961 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1962 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_981 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1962 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1961 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1963 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1964 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_982 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1964 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1963 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1965 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1966 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_983 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1966 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1965 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1967 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1968 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_984 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1968 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1967 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_246 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_984 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_983 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_982 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_981 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1969 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1970 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_985 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1970 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1969 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1971 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1972 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_986 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1972 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1971 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1973 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1974 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_987 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1974 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1973 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1975 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1976 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_988 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1976 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1975 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_247 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_988 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_987 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_986 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_985 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1977 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1978 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_989 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1978 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1977 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1979 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1980 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_990 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1980 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1979 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1981 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1982 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_991 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1982 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1981 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1983 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1984 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_992 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1984 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1983 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_248 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_992 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_991 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_990 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_989 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_62 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_248 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_247 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_246 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_245 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_1985 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1986 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_993 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1986 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1985 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1987 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1988 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_994 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1988 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1987 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1989 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1990 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_995 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1990 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1989 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1991 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_1992 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_996 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1992 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1991 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_249 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_996 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_995 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_994 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_993 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_1993 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1994 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_997 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1994 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1993 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1995 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1996 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_998 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1996 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1995 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1997 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_1998 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_999 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_1998 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1997 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_1999 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2000 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1000 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2000 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_1999 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_250 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1000 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_999 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_998 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_997 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2001 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2002 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1001 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2002 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2001 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2003 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2004 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1002 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2004 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2003 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2005 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2006 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1003 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2006 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2005 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2007 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2008 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1004 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2008 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2007 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_251 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1004 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1003 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1002 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1001 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2009 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2010 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1005 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2010 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2009 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2011 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2012 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1006 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2012 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2011 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2013 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2014 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1007 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2014 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2013 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2015 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2016 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1008 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2016 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2015 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_252 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1008 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1007 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1006 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1005 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_63 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_252 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_251 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_250 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_249 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_2017 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2018 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1009 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2018 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2017 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2019 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2020 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1010 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2020 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2019 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2021 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2022 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1011 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2022 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2021 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2023 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2024 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1012 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2024 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2023 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_253 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1012 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1011 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1010 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1009 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2025 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2026 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1013 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2026 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2025 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2027 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2028 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1014 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2028 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2027 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2029 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2030 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1015 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2030 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2029 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2031 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2032 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1016 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2032 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2031 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_254 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1016 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1015 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1014 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1013 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2033 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2034 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1017 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2034 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2033 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2035 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2036 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1018 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2036 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2035 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2037 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2038 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1019 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2038 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2037 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2039 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2040 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1020 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2040 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2039 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_255 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1020 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1019 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1018 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1017 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2041 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2042 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1021 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2042 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2041 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2043 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2044 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1022 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2044 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2043 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2045 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2046 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1023 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2046 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2045 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2047 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2048 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1024 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2048 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2047 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_256 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1024 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1023 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1022 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1021 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_64 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_256 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_255 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_254 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_253 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_16 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n4, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_64 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_63 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_62 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_61 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in8), .Z(n4) );
  CAOR2X1 U6 ( .A(s84[3]), .B(n5), .C(s83[3]), .D(n1), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n5), .C(s83[2]), .D(n1), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n5), .C(s83[1]), .D(n1), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n5), .C(s83[0]), .D(n1), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n4), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n4), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n4), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n4), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n5), .C(c_out810), .D(n1), .Z(c_out8) );
  CANR2X1 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n4), .Z(n1) );
endmodule


module bit32_4 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   n2, c1, c2, c3;

  bit8_16 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8(a32[7:0]), .b8(b32[7:0]), 
        .c_in8(c_in32) );
  bit8_15 A322 ( .sum8(sum32[15:8]), .c_out8(c2), .a8(a32[15:8]), .b8(
        b32[15:8]), .c_in8(c1) );
  bit8_14 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8(a32[23:16]), .b8(
        b32[23:16]), .c_in8(c2) );
  bit8_13 A324 ( .sum8({sum32[31:25], n2}), .c_out8(c_out32), .a8(a32[31:24]), 
        .b8(b32[31:24]), .c_in8(c3) );
  CNIVX4 U1 ( .A(n2), .Z(sum32[24]) );
endmodule


module Add_half_2049 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2050 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1025 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2050 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2049 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2051 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2052 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1026 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2052 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2051 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2053 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2054 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1027 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2054 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2053 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2055 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2056 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1028 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2056 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2055 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_257 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1028 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1027 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1026 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1025 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2057 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2058 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1029 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2058 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2057 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2059 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2060 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1030 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2060 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2059 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2061 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2062 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1031 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2062 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2061 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2063 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2064 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1032 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2064 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2063 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_258 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1032 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1031 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1030 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1029 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2065 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2066 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1033 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2066 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2065 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2067 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2068 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1034 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2068 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2067 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2069 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2070 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1035 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2070 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2069 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2071 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2072 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1036 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2072 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2071 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_259 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1036 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1035 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1034 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1033 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_2073 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2074 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1037 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2074 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2073 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2075 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2076 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1038 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2076 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2075 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2077 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2078 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1039 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2078 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2077 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2079 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2080 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1040 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2080 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2079 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_260 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1040 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1039 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1038 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1037 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n4) );
endmodule


module bit4_65 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_260 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_259 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_258 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_257 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CMX2X1 U4 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U7 ( .A(s43[0]), .Z(n3) );
  CIVX2 U8 ( .A(s44[0]), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n1), .Z(sum4[2]) );
  CIVX2 U10 ( .A(s43[1]), .Z(n5) );
  CIVX2 U11 ( .A(s44[1]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(n1), .Z(sum4[3]) );
endmodule


module Add_half_2081 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2082 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1041 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2082 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2081 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2083 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2084 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1042 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2084 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2083 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2085 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2086 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1043 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2086 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2085 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2087 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2088 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1044 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2088 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2087 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_261 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1044 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1043 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1042 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1041 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2089 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2090 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1045 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2090 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2089 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2091 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2092 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1046 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2092 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2091 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2093 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2094 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1047 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2094 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2093 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2095 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2096 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1048 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2096 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2095 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_262 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1048 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1047 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1046 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1045 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2097 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2098 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1049 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2098 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2097 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2099 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2100 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1050 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2100 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2099 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2101 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2102 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1051 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2102 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2101 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2103 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2104 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1052 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2104 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2103 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_263 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1052 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1051 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1050 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1049 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2105 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2106 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1053 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2106 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2105 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2107 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2108 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1054 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2108 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2107 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2109 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2110 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1055 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2110 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2109 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2111 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2112 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1056 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2112 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2111 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_264 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_1056 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1055 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1054 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1053 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
endmodule


module bit4_66 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_264 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_263 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_262 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_261 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CMX2X1 U5 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(s41[0]), .Z(n3) );
  CIVX2 U8 ( .A(s42[0]), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U10 ( .A(s41[1]), .Z(n5) );
  CIVX2 U11 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
endmodule


module Add_half_2113 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2114 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1057 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2114 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2113 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2115 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2116 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1058 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2116 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2115 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2117 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2118 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1059 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2118 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2117 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2119 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2120 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1060 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2120 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2119 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_265 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1060 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1059 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1058 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1057 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U7 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_2121 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2122 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1061 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2122 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2121 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2123 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2124 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1062 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2124 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2123 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2125 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2126 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1063 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2126 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2125 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2127 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2128 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1064 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2128 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2127 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_266 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1064 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1063 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1062 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1061 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_2129 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2130 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1065 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2130 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2129 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2131 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2132 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1066 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2132 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2131 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2133 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(n2) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U4 ( .A(b), .B(n2), .Z(sum) );
endmodule


module Add_half_2134 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1067 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2134 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2133 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2135 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(n1), .Z(sum) );
endmodule


module Add_half_2136 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1068 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2136 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2135 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_267 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1068 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1067 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1066 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1065 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
  CIVX1 U4 ( .A(n1), .Z(n6) );
  CIVX1 U5 ( .A(s2), .Z(n4) );
  CIVX1 U6 ( .A(s1), .Z(n5) );
  CIVX2 U7 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s3), .Z(n8) );
  CIVX2 U13 ( .A(s4), .Z(n7) );
endmodule


module Add_half_2137 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2138 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1069 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2138 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2137 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2139 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2140 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1070 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2140 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2139 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2141 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2142 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1071 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2142 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2141 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2143 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2144 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1072 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2144 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2143 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_268 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1072 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1071 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1070 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1069 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_67 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_268 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_267 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_266 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_265 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out4) );
  CIVX1 U4 ( .A(n1), .Z(n6) );
  CMX2XL U5 ( .A0(s43[1]), .A1(s44[1]), .S(n6), .Z(sum4[3]) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U7 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U8 ( .A(c_out410), .Z(n3) );
  CIVX2 U9 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U11 ( .A(s43[0]), .Z(n5) );
  CIVX2 U12 ( .A(s44[0]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(n6), .Z(sum4[2]) );
endmodule


module Add_half_2145 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2146 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1073 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2146 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2145 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2147 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2148 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1074 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2148 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2147 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2149 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2150 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1075 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2150 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2149 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2151 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2152 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1076 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2152 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2151 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_269 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1076 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1075 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1074 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1073 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CIVX2 U7 ( .A(s1), .Z(n3) );
  CIVX2 U8 ( .A(s2), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_2153 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2154 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1077 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2154 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2153 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2155 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2156 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1078 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2156 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2155 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2157 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2158 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1079 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2158 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2157 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2159 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2160 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1080 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2160 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2159 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_270 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1080 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1079 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1078 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1077 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_2161 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2162 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1081 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2162 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2161 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2163 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2164 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1082 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2164 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2163 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2165 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2166 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1083 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2166 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2165 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2167 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2168 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1084 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2168 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2167 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_271 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1084 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1083 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1082 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1081 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2169 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2170 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1085 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2170 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2169 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2171 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2172 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1086 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2172 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2171 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2173 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2174 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1087 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2174 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2173 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2175 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2176 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1088 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2176 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2175 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_272 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1088 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1087 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1086 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1085 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX1 U5 ( .A(n1), .Z(n4) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_68 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_272 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_271 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_270 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_269 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(n2), .Z(n1) );
  CIVX1 U4 ( .A(s41[0]), .Z(n6) );
  CMXI2X1 U5 ( .A0(n4), .A1(n3), .S(n1), .Z(c_out4) );
  CIVX2 U6 ( .A(c_out410), .Z(n4) );
  CIVX2 U7 ( .A(c_out411), .Z(n3) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CIVX2 U9 ( .A(s42[0]), .Z(n5) );
  CMXI2X1 U10 ( .A0(n6), .A1(n5), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U11 ( .A(s41[1]), .Z(n8) );
  CIVX2 U12 ( .A(s42[1]), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n10) );
  CIVX2 U15 ( .A(s44[0]), .Z(n9) );
  CMXI2X1 U16 ( .A0(n10), .A1(n9), .S(n1), .Z(sum4[2]) );
  CIVX2 U17 ( .A(s43[1]), .Z(n12) );
  CIVX2 U18 ( .A(s44[1]), .Z(n11) );
  CMXI2X1 U19 ( .A0(n12), .A1(n11), .S(n1), .Z(sum4[3]) );
endmodule


module bit8_17 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   n9, c_out800, c_out801, c_out810, c_out811, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_68 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_67 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_66 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_65 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X2 U3 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2X2 U4 ( .A0(s83[0]), .A1(s84[0]), .S(n2), .Z(sum8[4]) );
  CMXI2XL U5 ( .A0(n4), .A1(n3), .S(n2), .Z(c_out8) );
  CMX2X1 U6 ( .A0(s83[2]), .A1(s84[2]), .S(n2), .Z(sum8[6]) );
  CMXI2X1 U7 ( .A0(n8), .A1(n7), .S(c_in8), .Z(sum8[2]) );
  CIVX1 U8 ( .A(s81[2]), .Z(n8) );
  CIVX1 U9 ( .A(s82[2]), .Z(n7) );
  CMX2X2 U10 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n2) );
  CNIVX4 U11 ( .A(n9), .Z(sum8[0]) );
  CMXI2X1 U12 ( .A0(n6), .A1(n5), .S(c_in8), .Z(n9) );
  CMX2X1 U13 ( .A0(s83[3]), .A1(s84[3]), .S(n2), .Z(sum8[7]) );
  CMX2X1 U14 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2X1 U15 ( .A0(s83[1]), .A1(s84[1]), .S(n2), .Z(sum8[5]) );
  CIVX2 U16 ( .A(c_out810), .Z(n4) );
  CIVX2 U17 ( .A(c_out811), .Z(n3) );
  CIVX2 U18 ( .A(s81[0]), .Z(n6) );
  CIVX2 U19 ( .A(s82[0]), .Z(n5) );
endmodule


module Add_half_2177 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2178 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1089 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2178 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2177 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2179 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2180 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1090 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2180 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2179 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2181 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2182 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1091 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2182 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2181 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2183 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2184 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1092 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2184 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2183 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_273 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1092 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1091 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1090 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1089 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_2185 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2186 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1093 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2186 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2185 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2187 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2188 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1094 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2188 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2187 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2189 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2190 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1095 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2190 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2189 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2191 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2192 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1096 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2192 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2191 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_274 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1096 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1095 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1094 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1093 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_2193 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2194 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1097 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2194 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2193 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2195 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2196 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1098 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2196 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2195 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2197 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2198 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1099 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2198 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2197 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2199 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2200 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1100 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2200 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2199 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_275 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1100 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1099 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1098 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1097 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U4 ( .A(n1), .Z(n6) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_2201 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2202 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1101 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2202 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2201 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2203 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2204 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1102 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2204 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2203 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2205 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2206 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1103 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2206 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2205 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2207 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2208 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1104 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2208 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2207 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_276 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1104 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1103 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1102 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1101 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n4) );
endmodule


module bit4_69 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_276 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_275 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_274 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_273 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMX2XL U4 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2XL U5 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U6 ( .A0(c_out410), .A1(c_out411), .S(n4), .Z(c_out4) );
  CMX2X1 U7 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CIVX2 U9 ( .A(s41[1]), .Z(n3) );
  CIVX2 U10 ( .A(s42[1]), .Z(n2) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(c_in4), .Z(sum4[1]) );
endmodule


module Add_half_2209 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2210 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1105 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2210 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2209 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2211 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2212 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1106 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2212 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2211 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2213 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2214 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1107 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2214 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2213 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2215 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2216 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1108 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2216 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2215 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_277 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1108 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1107 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1106 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1105 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_2217 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2218 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1109 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2218 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2217 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2219 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2220 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1110 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2220 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2219 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2221 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2222 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1111 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2222 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2221 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2223 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2224 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1112 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2224 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2223 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_278 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1112 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1111 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1110 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1109 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_2225 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2226 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1113 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2226 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2225 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2227 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2228 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1114 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2228 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2227 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2229 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2230 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1115 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2230 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2229 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_2231 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2232 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1116 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2232 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2231 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_279 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1116 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1115 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1114 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1113 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n4) );
  CMXI2XL U4 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module Add_half_2233 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2234 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1117 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2234 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2233 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2235 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2236 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1118 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2236 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2235 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2237 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2238 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1119 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2238 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2237 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2239 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2240 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1120 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2240 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2239 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_280 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1120 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1119 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1118 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1117 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_70 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_280 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_279 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_278 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_277 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
  CIVX1 U4 ( .A(s41[0]), .Z(n5) );
  CIVX1 U5 ( .A(s42[0]), .Z(n4) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n8) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U13 ( .A(s43[0]), .Z(n7) );
  CIVX2 U14 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U15 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX2 U16 ( .A(s43[1]), .Z(n10) );
  CIVX2 U17 ( .A(s44[1]), .Z(n9) );
endmodule


module Add_half_2241 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2242 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1121 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2242 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2241 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2243 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2244 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1122 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2244 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2243 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2245 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2246 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1123 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2246 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2245 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2247 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2248 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1124 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2248 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2247 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_281 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1124 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1123 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1122 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1121 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2XL U4 ( .A0(n7), .A1(n6), .S(n1), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n7) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
endmodule


module Add_half_2249 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2250 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1125 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2250 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2249 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2251 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2252 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1126 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2252 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2251 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2253 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2254 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1127 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2254 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2253 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2255 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2256 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1128 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2256 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2255 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_282 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_1128 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1127 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1126 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1125 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
endmodule


module Add_half_2257 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2258 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1129 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2258 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2257 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2259 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2260 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1130 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2260 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2259 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2261 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2262 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1131 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2262 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2261 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2263 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2264 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1132 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2264 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2263 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_283 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1132 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1131 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1130 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1129 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s2), .Z(n4) );
  CIVX1 U4 ( .A(s1), .Z(n5) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n6) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_2265 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2266 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1133 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2266 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2265 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2267 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2268 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1134 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2268 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2267 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2269 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2270 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1135 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2270 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2269 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2271 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2272 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1136 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2272 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2271 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_284 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1136 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1135 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1134 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1133 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n4) );
  CIVX2 U8 ( .A(c_out11), .Z(n3) );
  CIVX2 U9 ( .A(n2), .Z(n5) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(n5), .Z(c_out2) );
endmodule


module bit4_71 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_284 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_283 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_282 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_281 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n6) );
  CIVX1 U4 ( .A(c_out411), .Z(n2) );
  CMX2XL U5 ( .A0(s43[1]), .A1(s44[1]), .S(n6), .Z(sum4[3]) );
  CMX2XL U6 ( .A0(s43[0]), .A1(s44[0]), .S(n6), .Z(sum4[2]) );
  CMX2X1 U7 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U8 ( .A(c_out410), .Z(n3) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out4) );
  CIVX2 U11 ( .A(s41[1]), .Z(n5) );
  CIVX2 U12 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
endmodule


module Add_half_2273 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2274 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1137 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2274 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2273 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2275 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2276 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1138 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2276 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2275 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2277 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2278 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1139 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2278 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2277 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2279 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2280 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1140 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2280 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2279 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_285 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1140 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1139 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1138 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1137 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2281 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2282 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1141 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2282 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2281 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2283 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2284 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1142 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2284 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2283 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2285 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2286 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1143 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2286 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2285 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2287 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2288 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1144 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2288 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2287 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_286 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1144 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1143 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1142 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1141 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2289 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2290 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1145 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2290 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2289 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2291 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2292 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1146 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2292 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2291 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2293 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2294 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1147 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2294 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2293 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2295 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2296 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1148 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2296 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2295 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_287 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1148 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1147 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1146 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1145 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n5), .A1(n6), .S(n1), .Z(sum2[1]) );
  CIVX1 U4 ( .A(n1), .Z(n4) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module Add_half_2297 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2298 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1149 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2298 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2297 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2299 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2300 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1150 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2300 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2299 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2301 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2302 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1151 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2302 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2301 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2303 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2304 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1152 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2304 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2303 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_288 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1152 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1151 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1150 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1149 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX1 U5 ( .A(n1), .Z(n4) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_72 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_288 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_287 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_286 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_285 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CMXI2XL U4 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n8) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U11 ( .A(s41[0]), .Z(n5) );
  CIVX2 U12 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n7) );
  CIVX2 U15 ( .A(s44[0]), .Z(n6) );
  CIVX2 U16 ( .A(s43[1]), .Z(n10) );
  CIVX2 U17 ( .A(s44[1]), .Z(n9) );
endmodule


module bit8_18 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_72 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4({b8[3], n5, 
        b8[1:0]}), .c_in4(1'b0) );
  bit4_71 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4({b8[3], n5, 
        b8[1:0]}), .c_in4(1'b1) );
  bit4_70 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_69 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X2 U3 ( .A0(s83[2]), .A1(s84[2]), .S(n6), .Z(sum8[6]) );
  CIVDXL U4 ( .A(c_in8), .Z0(n2), .Z1(n3) );
  CMX2X2 U5 ( .A0(s82[2]), .A1(s81[2]), .S(n2), .Z(sum8[2]) );
  CIVX2 U6 ( .A(b8[2]), .Z(n4) );
  CIVX4 U7 ( .A(n4), .Z(n5) );
  CMX2X1 U8 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n6) );
  CMXI2X1 U9 ( .A0(n9), .A1(n8), .S(c_in8), .Z(sum8[0]) );
  CMX2X2 U10 ( .A0(s83[1]), .A1(s84[1]), .S(n6), .Z(sum8[5]) );
  CIVX2 U11 ( .A(n7), .Z(n12) );
  CMXI2X1 U12 ( .A0(n11), .A1(n10), .S(n12), .Z(sum8[4]) );
  CMX2X2 U13 ( .A0(c_out810), .A1(c_out811), .S(n12), .Z(c_out8) );
  CMX2X1 U14 ( .A0(s83[3]), .A1(s84[3]), .S(n6), .Z(sum8[7]) );
  CMX2X1 U15 ( .A0(s81[3]), .A1(s82[3]), .S(n3), .Z(sum8[3]) );
  CMX2X1 U16 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMXI2X1 U17 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n7) );
  CIVX2 U18 ( .A(s81[0]), .Z(n9) );
  CIVX2 U19 ( .A(s82[0]), .Z(n8) );
  CIVX2 U20 ( .A(s83[0]), .Z(n11) );
  CIVX2 U21 ( .A(s84[0]), .Z(n10) );
endmodule


module Add_half_2305 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2306 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1153 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2306 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2305 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2307 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2308 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1154 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2308 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2307 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2309 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2310 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1155 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2310 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2309 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2311 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2312 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1156 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2312 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2311 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_289 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1156 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1155 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1154 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1153 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2313 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2314 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1157 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2314 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2313 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2315 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2316 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1158 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2316 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2315 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2317 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2318 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1159 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2318 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2317 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2319 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2320 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1160 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2320 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2319 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_290 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1160 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1159 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1158 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1157 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n2) );
  CMX2XL U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_2321 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2322 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1161 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2322 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2321 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2323 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2324 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1162 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2324 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2323 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2325 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2326 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1163 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2326 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2325 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2327 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2328 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1164 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2328 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2327 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_291 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1164 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1163 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1162 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1161 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n6) );
  CIVX1 U4 ( .A(s2), .Z(n4) );
  CIVX1 U5 ( .A(s1), .Z(n5) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U7 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_2329 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2330 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1165 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2330 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2329 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2331 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2332 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1166 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2332 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2331 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2333 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2334 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1167 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2334 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2333 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2335 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOX1 U1 ( .A(n1), .B(b), .Z(sum) );
  CNIVX1 U2 ( .A(a), .Z(n1) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2336 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1168 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2336 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2335 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_292 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1168 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1167 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1166 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1165 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_73 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_292 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_291 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_290 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_289 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CNIVX1 U3 ( .A(n2), .Z(n1) );
  CIVX1 U4 ( .A(n3), .Z(n2) );
  CMXI2X1 U5 ( .A0(n7), .A1(n6), .S(n1), .Z(sum4[2]) );
  CMXI2XL U6 ( .A0(n9), .A1(n8), .S(n1), .Z(sum4[3]) );
  CMX2X1 U7 ( .A0(c_out410), .A1(c_out411), .S(n2), .Z(c_out4) );
  CMX2X1 U8 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX1 U9 ( .A(s43[1]), .Z(n9) );
  CMXI2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n3) );
  CIVX2 U11 ( .A(s41[1]), .Z(n5) );
  CIVX2 U12 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n7) );
  CIVX2 U15 ( .A(s44[0]), .Z(n6) );
  CIVX2 U16 ( .A(s44[1]), .Z(n8) );
endmodule


module Add_half_2337 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2338 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1169 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2338 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2337 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2339 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2340 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1170 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2340 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2339 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2341 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2342 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1171 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2342 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2341 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2343 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2344 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1172 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2344 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2343 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_293 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1172 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1171 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1170 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1169 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_2345 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2346 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1173 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2346 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2345 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2347 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2348 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1174 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2348 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2347 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2349 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2350 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1175 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2350 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2349 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2351 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2352 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1176 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2352 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2351 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_294 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1176 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1175 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1174 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1173 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2353 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2354 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1177 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2354 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2353 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2355 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2356 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1178 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2356 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2355 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2357 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2358 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1179 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2358 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2357 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2359 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2360 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1180 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2360 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2359 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_295 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n2, n3, n4, n5,
         n6, n7;

  Add_full_1180 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1179 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1178 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1177 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CIVDXL U4 ( .A(n2), .Z0(n5) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n4) );
  CIVX2 U7 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX2 U9 ( .A(s3), .Z(n7) );
  CIVX2 U10 ( .A(s4), .Z(n6) );
  CMXI2X1 U11 ( .A0(n7), .A1(n6), .S(n5), .Z(sum2[1]) );
endmodule


module Add_half_2361 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2362 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1181 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2362 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2361 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2363 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2364 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1182 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2364 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2363 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2365 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2366 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1183 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2366 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2365 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2367 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2368 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1184 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2368 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2367 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_296 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1184 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1183 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1182 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1181 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_74 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_296 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_295 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_294 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_293 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2X1 U4 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out4) );
  CMX2XL U5 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U6 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2X1 U7 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U8 ( .A(c_out410), .Z(n4) );
  CIVX2 U9 ( .A(c_out411), .Z(n3) );
  CMXI2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CIVX2 U11 ( .A(s41[0]), .Z(n6) );
  CIVX2 U12 ( .A(s42[0]), .Z(n5) );
  CMXI2X1 U13 ( .A0(n6), .A1(n5), .S(c_in4), .Z(sum4[0]) );
endmodule


module Add_half_2369 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2370 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1185 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2370 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2369 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2371 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2372 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1186 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2372 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2371 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2373 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2374 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1187 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2374 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2373 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2375 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2376 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1188 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2376 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2375 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_297 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1188 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1187 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1186 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1185 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CIVX2 U7 ( .A(s1), .Z(n3) );
  CIVX2 U8 ( .A(s2), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module Add_half_2377 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2378 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1189 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2378 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2377 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2379 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2380 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1190 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2380 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2379 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2381 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2382 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1191 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2382 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2381 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2383 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2384 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1192 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2384 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2383 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_298 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1192 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1191 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1190 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1189 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_2385 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2386 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1193 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2386 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2385 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2387 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2388 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1194 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2388 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2387 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2389 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2390 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1195 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2390 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2389 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2391 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2392 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1196 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2392 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2391 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_299 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1196 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1195 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1194 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1193 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_2393 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2394 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1197 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2394 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2393 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2395 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2396 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1198 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2396 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2395 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2397 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2398 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1199 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2398 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2397 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2399 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2400 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1200 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2400 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2399 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_300 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1200 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1199 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1198 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1197 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_75 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_300 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_299 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_298 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_297 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n6), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n6), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n6) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out4) );
  CIVX2 U11 ( .A(s41[0]), .Z(n5) );
  CIVX2 U12 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
endmodule


module Add_half_2401 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2402 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1201 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2402 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2401 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2403 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2404 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1202 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2404 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2403 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2405 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2406 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1203 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2406 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2405 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_2407 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2408 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1204 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2408 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2407 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_301 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1204 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1203 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1202 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1201 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_2409 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2410 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1205 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2410 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2409 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2411 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2412 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1206 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2412 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2411 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2413 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2414 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1207 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2414 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2413 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2415 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2416 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2, n3;

  CEOX1 U1 ( .A(a), .B(n3), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(n3), .Z(c_out) );
  CIVXL U3 ( .A(b), .Z(n2) );
  CIVX2 U4 ( .A(n2), .Z(n3) );
endmodule


module Add_full_1208 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2416 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2415 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_302 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1208 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1207 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1206 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1205 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(n1), .Z(n2) );
  CMX2X1 U4 ( .A0(c_out11), .A1(c_out10), .S(n1), .Z(c_out2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_2417 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2418 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1209 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2418 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2417 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2419 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2420 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1210 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2420 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2419 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2421 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2422 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1211 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2422 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2421 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2423 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2424 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1212 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2424 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2423 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_303 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1212 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1211 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1210 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1209 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2425 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2426 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1213 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2426 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2425 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2427 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2428 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1214 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2428 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2427 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2429 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2430 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1215 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2430 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2429 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2431 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2432 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1216 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2432 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2431 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_304 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1216 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1215 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1214 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1213 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module bit4_76 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_304 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_303 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_302 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_301 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n8), .Z(sum4[3]) );
  CMX2X1 U4 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U5 ( .A(c_out410), .Z(n3) );
  CIVX2 U6 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n8) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U10 ( .A(s41[1]), .Z(n5) );
  CIVX2 U11 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U13 ( .A(s43[0]), .Z(n7) );
  CIVX2 U14 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U15 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
endmodule


module bit8_19 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_76 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_75 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_74 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_73 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X1 U3 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CMX2X2 U4 ( .A0(s83[1]), .A1(s84[1]), .S(n1), .Z(sum8[5]) );
  CMXI2X1 U5 ( .A0(c_out810), .A1(c_out811), .S(n4), .Z(n2) );
  CIVX2 U6 ( .A(n2), .Z(c_out8) );
  CMXI2X1 U7 ( .A0(s83[0]), .A1(s84[0]), .S(n4), .Z(n3) );
  CIVX3 U8 ( .A(n3), .Z(sum8[4]) );
  CIVX1 U9 ( .A(s84[2]), .Z(n7) );
  CIVX1 U10 ( .A(s83[2]), .Z(n8) );
  CMXI2X2 U11 ( .A0(n8), .A1(n7), .S(n1), .Z(sum8[6]) );
  CMX2X2 U12 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n4) );
  CMX2X2 U13 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2X2 U14 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2X2 U15 ( .A0(s81[0]), .A1(s82[0]), .S(c_in8), .Z(sum8[0]) );
  CMX2X1 U16 ( .A0(s83[3]), .A1(s84[3]), .S(n1), .Z(sum8[7]) );
  CIVX2 U17 ( .A(s81[3]), .Z(n6) );
  CIVX2 U18 ( .A(s82[3]), .Z(n5) );
  CMXI2X1 U19 ( .A0(n6), .A1(n5), .S(c_in8), .Z(sum8[3]) );
endmodule


module Add_half_2433 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2434 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1217 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2434 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2433 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2435 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2436 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1218 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2436 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2435 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2437 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2438 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1219 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2438 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2437 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2439 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2440 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1220 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2440 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2439 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_305 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1220 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1219 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1218 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1217 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2441 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2442 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1221 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2442 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2441 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2443 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2444 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1222 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2444 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2443 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2445 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2446 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1223 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2446 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2445 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2447 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2448 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1224 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2448 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2447 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_306 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1224 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1223 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1222 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1221 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2449 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2450 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1225 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2450 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2449 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2451 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2452 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1226 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2452 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2451 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2453 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2454 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1227 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2454 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2453 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2455 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2456 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1228 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2456 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2455 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_307 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1228 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1227 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1226 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1225 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2457 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2458 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1229 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2458 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2457 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2459 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2460 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1230 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2460 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2459 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2461 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2462 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1231 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2462 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2461 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2463 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2464 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1232 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2464 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2463 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_308 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1232 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1231 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1230 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1229 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_77 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_308 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_307 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_306 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_305 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_2465 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2466 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1233 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2466 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2465 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2467 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2468 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1234 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2468 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2467 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2469 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2470 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1235 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2470 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2469 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2471 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2472 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1236 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2472 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2471 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_309 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1236 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1235 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1234 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1233 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2473 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2474 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1237 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2474 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2473 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2475 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2476 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1238 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2476 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2475 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2477 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2478 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1239 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2478 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2477 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2479 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2480 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1240 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2480 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2479 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_310 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1240 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1239 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1238 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1237 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2481 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2482 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1241 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2482 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2481 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2483 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2484 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1242 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2484 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2483 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2485 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2486 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1243 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2486 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2485 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2487 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2488 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1244 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2488 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2487 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_311 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1244 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1243 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1242 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1241 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2489 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2490 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1245 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2490 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2489 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2491 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2492 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1246 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2492 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2491 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2493 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2494 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1247 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2494 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2493 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2495 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2496 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1248 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2496 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2495 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_312 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1248 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1247 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1246 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1245 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_78 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_312 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_311 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_310 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_309 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_2497 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2498 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1249 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2498 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2497 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2499 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2500 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1250 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2500 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2499 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2501 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2502 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1251 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2502 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2501 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2503 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2504 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1252 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2504 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2503 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_313 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1252 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1251 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1250 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1249 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2505 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2506 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1253 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2506 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2505 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2507 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2508 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1254 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2508 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2507 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2509 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2510 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1255 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2510 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2509 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2511 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2512 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1256 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2512 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2511 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_314 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1256 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1255 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1254 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1253 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2513 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2514 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1257 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2514 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2513 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2515 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2516 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1258 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2516 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2515 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2517 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2518 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1259 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2518 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2517 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2519 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2520 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1260 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2520 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2519 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_315 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1260 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1259 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1258 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1257 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2521 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2522 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1261 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2522 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2521 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2523 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2524 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1262 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2524 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2523 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2525 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2526 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1263 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2526 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2525 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2527 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2528 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1264 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2528 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2527 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_316 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1264 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1263 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1262 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1261 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_79 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_316 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_315 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_314 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_313 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_2529 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2530 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1265 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2530 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2529 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2531 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2532 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1266 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2532 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2531 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2533 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2534 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1267 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2534 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2533 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2535 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2536 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1268 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2536 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2535 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_317 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1268 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1267 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1266 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1265 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2537 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2538 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1269 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2538 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2537 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2539 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2540 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1270 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2540 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2539 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2541 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2542 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1271 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2542 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2541 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2543 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2544 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1272 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2544 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2543 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_318 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1272 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1271 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1270 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1269 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2545 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2546 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1273 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2546 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2545 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2547 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2548 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1274 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2548 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2547 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2549 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2550 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1275 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2550 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2549 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2551 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2552 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1276 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2552 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2551 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_319 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1276 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1275 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1274 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1273 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_2553 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2554 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1277 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2554 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2553 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2555 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2556 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1278 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2556 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2555 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2557 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2558 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1279 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2558 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2557 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2559 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2560 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1280 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2560 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2559 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_320 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1280 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1279 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1278 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1277 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_80 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_320 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_319 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_318 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_317 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_20 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n4, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_80 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_79 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_78 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_77 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in8), .Z(n4) );
  CAOR2X1 U6 ( .A(s84[3]), .B(n5), .C(s83[3]), .D(n1), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n5), .C(s83[2]), .D(n1), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n5), .C(s83[1]), .D(n1), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n5), .C(s83[0]), .D(n1), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n4), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n4), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n4), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n4), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n5), .C(c_out810), .D(n1), .Z(c_out8) );
  CANR2X1 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n4), .Z(n1) );
endmodule


module bit32_5 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   c1, c2, c3;

  bit8_20 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8(a32[7:0]), .b8(b32[7:0]), 
        .c_in8(c_in32) );
  bit8_19 A322 ( .sum8(sum32[15:8]), .c_out8(c2), .a8(a32[15:8]), .b8(
        b32[15:8]), .c_in8(c1) );
  bit8_18 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8(a32[23:16]), .b8(
        b32[23:16]), .c_in8(c2) );
  bit8_17 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8(a32[31:24]), .b8(
        b32[31:24]), .c_in8(c3) );
endmodule


module Add_half_2561 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2562 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1281 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2562 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2561 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2563 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2564 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1282 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2564 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2563 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2565 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2566 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1283 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2566 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2565 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2567 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2568 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1284 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2568 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2567 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_321 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1284 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1283 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1282 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1281 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CIVX2 U5 ( .A(s1), .Z(n3) );
  CIVX2 U6 ( .A(s2), .Z(n2) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(s3), .Z(n5) );
  CIVX2 U9 ( .A(s4), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
endmodule


module Add_half_2569 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2570 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1285 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2570 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2569 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2571 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2572 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1286 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2572 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2571 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2573 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2574 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1287 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2574 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2573 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2575 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2576 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1288 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2576 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2575 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_322 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_1288 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1287 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1286 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1285 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CIVX1 U5 ( .A(s3), .Z(n3) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(s4), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(sum2[1]) );
endmodule


module Add_half_2577 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2578 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1289 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2578 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2577 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2579 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2580 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1290 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2580 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2579 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2581 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2582 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1291 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2582 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2581 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2583 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2584 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1292 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2584 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2583 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_323 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1292 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1291 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1290 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1289 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n7), .A1(n8), .S(n1), .Z(sum2[1]) );
  CMXI2XL U4 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX1 U5 ( .A(n1), .Z(n6) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s3), .Z(n8) );
  CIVX2 U13 ( .A(s4), .Z(n7) );
endmodule


module Add_half_2585 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2586 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1293 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2586 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2585 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2587 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2588 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1294 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2588 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2587 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2589 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2590 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1295 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2590 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2589 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2591 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2592 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1296 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2592 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2591 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_324 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1296 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1295 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1294 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1293 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX1 U6 ( .A(n1), .Z(n4) );
  CIVX2 U7 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module bit4_81 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_324 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_323 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_322 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_321 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U7 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
endmodule


module Add_half_2593 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2594 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1297 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2594 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2593 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2595 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2596 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1298 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2596 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2595 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2597 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2598 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1299 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2598 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2597 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2599 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2600 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1300 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2600 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2599 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_325 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_1300 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1299 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1298 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1297 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(s3), .Z(n3) );
  CIVX2 U7 ( .A(s4), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(sum2[1]) );
endmodule


module Add_half_2601 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2602 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1301 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2602 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2601 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2603 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2604 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1302 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2604 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2603 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2605 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2606 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1303 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2606 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2605 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_2607 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2608 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1304 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2608 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2607 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_326 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_1304 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1303 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1302 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1301 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CIVX1 U5 ( .A(s3), .Z(n3) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(s4), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(sum2[1]) );
endmodule


module Add_half_2609 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2610 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1305 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2610 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2609 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2611 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2612 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1306 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2612 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2611 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2613 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2614 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1307 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2614 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2613 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2615 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2616 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1308 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2616 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2615 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_327 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1308 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1307 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1306 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1305 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2617 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2618 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1309 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2618 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2617 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2619 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2620 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1310 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2620 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2619 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2621 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2622 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1311 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2622 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2621 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2623 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2624 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1312 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2624 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2623 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_328 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1312 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1311 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1310 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1309 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n4) );
  CMXI2X1 U4 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module bit4_82 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_328 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_327 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_326 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_325 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CMX2XL U4 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U6 ( .A(s41[0]), .Z(n3) );
  CIVX2 U7 ( .A(s42[0]), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U9 ( .A(s41[1]), .Z(n5) );
  CIVX2 U10 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(s43[0]), .Z(n7) );
  CIVX2 U13 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n1), .Z(sum4[2]) );
endmodule


module Add_half_2625 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2626 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1313 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2626 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2625 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2627 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2628 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1314 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2628 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2627 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2629 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2630 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1315 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2630 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2629 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2631 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2632 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1316 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2632 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2631 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_329 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1316 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1315 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1314 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1313 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U7 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_2633 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2634 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1317 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2634 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2633 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2635 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2636 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1318 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2636 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2635 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2637 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2638 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1319 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2638 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2637 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2639 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2640 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1320 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2640 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2639 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_330 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1320 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1319 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1318 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1317 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_2641 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2642 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1321 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2642 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2641 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2643 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2644 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1322 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2644 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2643 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2645 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2646 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1323 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2646 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2645 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2647 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2648 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1324 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2648 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2647 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_331 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1324 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1323 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1322 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1321 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(c_out11), .Z(n2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2649 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2650 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1325 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2650 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2649 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2651 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2652 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1326 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2652 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2651 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2653 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2654 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1327 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2654 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2653 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2655 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2656 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1328 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2656 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2655 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_332 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1328 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1327 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1326 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1325 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CIVX2 U4 ( .A(n2), .Z(n5) );
  CIVX1 U5 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(c_out10), .Z(n4) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(n5), .Z(c_out2) );
endmodule


module bit4_83 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_332 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_331 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_330 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_329 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(c_in4), .Z(n1) );
  CIVX1 U4 ( .A(s41[0]), .Z(n6) );
  CIVX2 U5 ( .A(n2), .Z(n11) );
  CMXI2XL U6 ( .A0(n13), .A1(n12), .S(n11), .Z(sum4[3]) );
  CMXI2X1 U7 ( .A0(c_out401), .A1(c_out400), .S(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_out410), .Z(n4) );
  CIVX2 U9 ( .A(c_out411), .Z(n3) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(n11), .Z(c_out4) );
  CIVX2 U11 ( .A(s42[0]), .Z(n5) );
  CMXI2X1 U12 ( .A0(n6), .A1(n5), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U13 ( .A(s41[1]), .Z(n8) );
  CIVX2 U14 ( .A(s42[1]), .Z(n7) );
  CMXI2X1 U15 ( .A0(n8), .A1(n7), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U16 ( .A(s43[0]), .Z(n10) );
  CIVX2 U17 ( .A(s44[0]), .Z(n9) );
  CMXI2X1 U18 ( .A0(n10), .A1(n9), .S(n11), .Z(sum4[2]) );
  CIVX2 U19 ( .A(s43[1]), .Z(n13) );
  CIVX2 U20 ( .A(s44[1]), .Z(n12) );
endmodule


module Add_half_2657 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2658 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1329 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2658 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2657 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2659 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2660 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1330 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2660 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2659 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2661 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2662 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1331 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2662 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2661 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2663 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2664 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1332 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2664 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2663 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_333 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1332 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1331 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1330 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1329 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CIVX2 U7 ( .A(s1), .Z(n3) );
  CIVX2 U8 ( .A(s2), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_2665 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2666 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1333 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2666 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2665 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2667 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2668 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1334 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2668 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2667 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2669 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2670 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1335 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2670 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2669 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2671 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2672 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1336 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2672 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2671 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_334 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1336 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1335 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1334 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1333 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_2673 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2674 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1337 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2674 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2673 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2675 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2676 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1338 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2676 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2675 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2677 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2678 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1339 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2678 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2677 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2679 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2680 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1340 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2680 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2679 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_335 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1340 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1339 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1338 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1337 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(n1), .Z(n6) );
  CIVX1 U5 ( .A(s4), .Z(n7) );
  CIVX1 U6 ( .A(s3), .Z(n8) );
  CIVX1 U7 ( .A(s2), .Z(n4) );
  CIVX1 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(c_out10), .Z(n3) );
  CIVX2 U10 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U11 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U12 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_2681 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2682 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1341 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2682 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2681 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2683 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2684 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1342 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2684 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2683 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2685 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2686 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1343 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2686 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2685 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2687 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2688 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1344 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2688 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2687 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_336 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1344 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1343 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1342 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1341 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_84 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_336 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_335 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_334 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_333 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2X1 U4 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out4) );
  CMX2XL U5 ( .A0(s43[1]), .A1(s44[1]), .S(n6), .Z(sum4[3]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U7 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX1 U8 ( .A(c_out410), .Z(n3) );
  CIVX2 U9 ( .A(c_out411), .Z(n2) );
  CIVX2 U10 ( .A(n1), .Z(n6) );
  CIVX2 U11 ( .A(s43[0]), .Z(n5) );
  CIVX2 U12 ( .A(s44[0]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(n6), .Z(sum4[2]) );
endmodule


module bit8_21 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   n16, c_out800, c_out801, c_out810, c_out811, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_84 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4({b8[3:2], n6, 
        b8[0]}), .c_in4(1'b0) );
  bit4_83 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4({b8[3:2], n6, 
        b8[0]}), .c_in4(1'b1) );
  bit4_82 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_81 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CNIVX4 U3 ( .A(n16), .Z(sum8[0]) );
  CIVX2 U4 ( .A(n7), .Z(n4) );
  CMX2X1 U5 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMXI2X1 U6 ( .A0(n11), .A1(n10), .S(c_in8), .Z(n16) );
  CMXI2X1 U7 ( .A0(n15), .A1(n14), .S(n5), .Z(sum8[7]) );
  CND2X2 U8 ( .A(s83[0]), .B(n4), .Z(n2) );
  CMX2X2 U9 ( .A0(s83[1]), .A1(s84[1]), .S(n7), .Z(sum8[5]) );
  CND2X4 U10 ( .A(n2), .B(n3), .Z(sum8[4]) );
  CND2X1 U11 ( .A(s84[0]), .B(n7), .Z(n3) );
  CMX2X1 U12 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n7) );
  CIVX1 U13 ( .A(n4), .Z(n5) );
  CNIVX3 U14 ( .A(b8[1]), .Z(n6) );
  CMXI2X1 U15 ( .A0(n13), .A1(n12), .S(c_in8), .Z(sum8[3]) );
  CMX2X2 U16 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2X2 U17 ( .A0(s83[2]), .A1(s84[2]), .S(n5), .Z(sum8[6]) );
  CIVXL U18 ( .A(s82[3]), .Z(n12) );
  CMXI2XL U19 ( .A0(n9), .A1(n8), .S(n5), .Z(c_out8) );
  CIVX2 U20 ( .A(c_out810), .Z(n9) );
  CIVX2 U21 ( .A(c_out811), .Z(n8) );
  CIVX2 U22 ( .A(s81[0]), .Z(n11) );
  CIVX2 U23 ( .A(s82[0]), .Z(n10) );
  CIVX2 U24 ( .A(s81[3]), .Z(n13) );
  CIVX2 U25 ( .A(s83[3]), .Z(n15) );
  CIVX2 U26 ( .A(s84[3]), .Z(n14) );
endmodule


module Add_half_2689 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2690 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1345 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2690 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2689 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2691 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2692 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1346 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2692 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2691 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2693 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVX1 U1 ( .A(a), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(n2) );
  CAN2X1 U3 ( .A(n2), .B(b), .Z(c_out) );
  CEOX1 U4 ( .A(n2), .B(b), .Z(sum) );
endmodule


module Add_half_2694 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1347 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2694 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2693 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2695 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2696 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1348 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2696 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2695 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_337 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1348 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1347 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1346 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1345 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_2697 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2698 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1349 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2698 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2697 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2699 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2700 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1350 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2700 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2699 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2701 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2702 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1351 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2702 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2701 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2703 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2704 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1352 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2704 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2703 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_338 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1352 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1351 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1350 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1349 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX1 U4 ( .A(c_out11), .Z(n2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n3) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n4) );
endmodule


module Add_half_2705 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2706 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1353 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2706 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2705 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2707 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2708 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1354 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2708 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2707 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2709 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2710 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1355 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2710 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2709 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2711 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2712 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1356 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2712 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2711 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_339 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1356 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1355 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1354 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1353 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CIVX2 U5 ( .A(c_out10), .Z(n4) );
  CIVX2 U6 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX2 U8 ( .A(s1), .Z(n6) );
  CIVX2 U9 ( .A(s2), .Z(n5) );
  CMXI2X1 U10 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n1), .Z(sum2[1]) );
endmodule


module Add_half_2713 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(a), .B(n2), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2714 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1357 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2714 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2713 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2715 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2716 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1358 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2716 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2715 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2717 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2718 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1359 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2718 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2717 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2719 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2720 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1360 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2720 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2719 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_340 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1360 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1359 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1358 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1357 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n4) );
  CIVX2 U8 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module bit4_85 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_340 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_339 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_338 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_337 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U7 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CIVX2 U8 ( .A(c_out410), .Z(n3) );
  CIVX2 U9 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module Add_half_2721 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2722 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1361 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2722 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2721 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2723 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2724 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1362 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2724 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2723 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2725 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2726 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1363 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2726 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2725 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2727 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2728 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1364 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2728 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2727 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_341 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1364 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1363 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1362 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1361 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2729 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2730 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1365 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2730 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2729 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2731 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2732 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1366 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2732 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2731 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2733 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2734 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1367 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2734 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2733 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2735 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2736 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1368 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2736 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2735 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_342 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1368 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1367 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1366 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1365 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2737 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2738 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1369 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2738 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2737 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2739 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2740 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1370 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2740 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2739 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2741 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2742 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1371 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2742 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2741 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2743 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2744 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1372 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2744 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2743 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_343 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1372 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1371 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1370 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1369 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2745 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2746 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1373 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2746 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2745 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2747 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2748 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1374 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2748 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2747 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2749 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2750 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1375 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2750 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2749 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2751 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2752 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n3), .B(n4), .Z(sum) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CND2XL U3 ( .A(n1), .B(b), .Z(n4) );
  CIVXL U4 ( .A(b), .Z(n2) );
  CIVXL U5 ( .A(a), .Z(n1) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1376 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2752 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2751 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_344 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1376 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1375 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1374 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1373 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_86 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_344 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_343 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_342 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_341 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(s41[1]), .Z(n7) );
  CMXI2XL U4 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(s43[0]), .A1(s44[0]), .S(n8), .Z(sum4[2]) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n8) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U11 ( .A(s41[0]), .Z(n5) );
  CIVX2 U12 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U14 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U15 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U16 ( .A(s43[1]), .Z(n10) );
  CIVX2 U17 ( .A(s44[1]), .Z(n9) );
endmodule


module Add_half_2753 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2754 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1377 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2754 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2753 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2755 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2756 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1378 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2756 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2755 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2757 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2758 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1379 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2758 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2757 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2759 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2760 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1380 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2760 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2759 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_345 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1380 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1379 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1378 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1377 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(n1), .Z(n4) );
  CIVX2 U6 ( .A(s1), .Z(n3) );
  CIVX2 U7 ( .A(s2), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_2761 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2762 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1381 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2762 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2761 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2763 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2764 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1382 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2764 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2763 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2765 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2766 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1383 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2766 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2765 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2767 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2768 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1384 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2768 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2767 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_346 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1384 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1383 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1382 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1381 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U7 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_2769 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2770 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1385 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2770 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2769 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2771 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2772 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1386 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2772 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2771 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2773 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2774 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVXL U1 ( .A(a), .Z(n1) );
  CND2X1 U2 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U3 ( .A(b), .Z(n2) );
  CND2XL U4 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U5 ( .A(a), .B(n2), .Z(n3) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1387 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2774 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2773 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2775 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2776 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1388 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2776 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2775 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CND2X1 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_347 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1388 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1387 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1386 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1385 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(n1), .Z(n6) );
  CIVX1 U4 ( .A(s1), .Z(n5) );
  CMXI2X1 U5 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_2777 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2778 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1389 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2778 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2777 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2779 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2780 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1390 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2780 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2779 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2781 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2782 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1391 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2782 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2781 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2783 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2784 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1392 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2784 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2783 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_348 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1392 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1391 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1390 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1389 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2X1 U3 ( .A(c_out10), .B(n1), .Z(n2) );
  CND2X1 U4 ( .A(c_out11), .B(n5), .Z(n3) );
  CND2X1 U5 ( .A(n2), .B(n3), .Z(c_out2) );
  CIVX1 U6 ( .A(n5), .Z(n1) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n4) );
  CIVX2 U10 ( .A(n4), .Z(n5) );
endmodule


module bit4_87 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_348 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_347 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_346 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_345 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMX2X1 U4 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2XL U5 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U7 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CIVX2 U9 ( .A(c_out410), .Z(n4) );
  CIVX2 U10 ( .A(c_out411), .Z(n3) );
  CMXI2X1 U11 ( .A0(n4), .A1(n3), .S(n2), .Z(c_out4) );
endmodule


module Add_half_2785 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2786 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1393 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2786 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2785 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2787 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2788 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1394 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2788 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2787 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2789 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2790 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1395 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2790 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2789 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_2791 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2792 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1396 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2792 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2791 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_349 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1396 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1395 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1394 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1393 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_2793 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2794 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1397 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2794 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2793 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2795 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2796 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1398 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2796 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2795 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2797 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2798 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1399 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2798 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2797 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_2799 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2800 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1400 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2800 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2799 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_350 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1400 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1399 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1398 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1397 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2801 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2802 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1401 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2802 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2801 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2803 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2804 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1402 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2804 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2803 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2805 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2806 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1403 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2806 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2805 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CND2X1 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_2807 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2808 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1404 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2808 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2807 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX1 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_351 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1404 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1403 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1402 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1401 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2809 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2810 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1405 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2810 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2809 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2811 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2812 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1406 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2812 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2811 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2813 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2814 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1407 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2814 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2813 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX1 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_2815 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2816 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n3), .B(n4), .Z(sum) );
  CND2XL U2 ( .A(n1), .B(b), .Z(n4) );
  CND2XL U3 ( .A(a), .B(n2), .Z(n3) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1408 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2816 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2815 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_352 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1408 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1407 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1406 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1405 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_88 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_352 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_351 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_350 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_349 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(s42[0]), .Z(n4) );
  CIVXL U4 ( .A(n1), .Z(n10) );
  CMXI2X1 U5 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out4) );
  CMXI2X1 U6 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CIVX1 U7 ( .A(c_out410), .Z(n3) );
  CIVX1 U8 ( .A(c_out411), .Z(n2) );
  CMXI2XL U9 ( .A0(n12), .A1(n11), .S(n10), .Z(sum4[3]) );
  CMXI2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U11 ( .A(s41[0]), .Z(n5) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U13 ( .A(s41[1]), .Z(n7) );
  CIVX2 U14 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U15 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U16 ( .A(s43[0]), .Z(n9) );
  CIVX2 U17 ( .A(s44[0]), .Z(n8) );
  CIVX2 U18 ( .A(s43[1]), .Z(n12) );
  CIVX2 U19 ( .A(s44[1]), .Z(n11) );
endmodule


module bit8_22 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_88 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_87 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_86 A83 ( .sum4(s83), .c_out4(c_out810), .a4({a8[7:5], n2}), .b4({n1, 
        b8[6:4]}), .c_in4(1'b0) );
  bit4_85 A84 ( .sum4(s84), .c_out4(c_out811), .a4({a8[7:5], n2}), .b4({n1, 
        b8[6:4]}), .c_in4(1'b1) );
  CND2X1 U3 ( .A(c_out811), .B(n15), .Z(n8) );
  CND2X2 U4 ( .A(s83[0]), .B(n6), .Z(n3) );
  CNIVX4 U5 ( .A(b8[7]), .Z(n1) );
  CND2X2 U6 ( .A(n7), .B(n8), .Z(c_out8) );
  CNIVX4 U7 ( .A(a8[4]), .Z(n2) );
  CMX2X2 U8 ( .A0(s81[3]), .A1(s82[3]), .S(n5), .Z(sum8[3]) );
  CMX2X2 U9 ( .A0(s83[3]), .A1(s84[3]), .S(n9), .Z(sum8[7]) );
  CMXI2X4 U10 ( .A0(n14), .A1(n13), .S(n15), .Z(sum8[5]) );
  CIVX2 U11 ( .A(n15), .Z(n6) );
  CMX2X2 U12 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CNIVX1 U13 ( .A(c_in8), .Z(n5) );
  CMX2X2 U14 ( .A0(s81[2]), .A1(s82[2]), .S(n5), .Z(sum8[2]) );
  CIVX1 U15 ( .A(s83[1]), .Z(n14) );
  CND2X1 U16 ( .A(s84[0]), .B(n15), .Z(n4) );
  CND2X4 U17 ( .A(n3), .B(n4), .Z(sum8[4]) );
  CMX2X2 U18 ( .A0(s83[2]), .A1(s84[2]), .S(n15), .Z(sum8[6]) );
  CND2X1 U19 ( .A(c_out810), .B(n6), .Z(n7) );
  CIVX2 U20 ( .A(n10), .Z(n15) );
  CIVXL U21 ( .A(n6), .Z(n9) );
  CMXI2X1 U22 ( .A0(n12), .A1(n11), .S(c_in8), .Z(sum8[0]) );
  CMXI2X1 U23 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n10) );
  CIVX2 U24 ( .A(s81[0]), .Z(n12) );
  CIVX2 U25 ( .A(s82[0]), .Z(n11) );
  CIVX2 U26 ( .A(s84[1]), .Z(n13) );
endmodule


module Add_half_2817 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2818 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1409 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2818 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2817 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2819 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2820 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1410 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2820 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2819 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2821 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2822 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1411 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2822 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2821 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2823 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2824 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1412 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2824 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2823 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_353 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1412 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1411 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1410 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1409 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_2825 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2826 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1413 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2826 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2825 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2827 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2828 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1414 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2828 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2827 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2829 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2830 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1415 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2830 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2829 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2831 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2832 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1416 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2832 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2831 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_354 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1416 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1415 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1414 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1413 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_2833 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2834 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1417 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2834 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2833 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2835 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2836 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1418 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2836 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2835 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2837 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2838 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1419 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2838 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2837 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2839 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2840 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1420 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2840 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2839 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_355 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1420 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1419 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1418 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1417 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CIVX1 U5 ( .A(s1), .Z(n6) );
  CIVXL U6 ( .A(n2), .Z(n7) );
  CMXI2X1 U7 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMX2XL U8 ( .A0(s3), .A1(s4), .S(n7), .Z(sum2[1]) );
  CIVX2 U9 ( .A(c_out10), .Z(n4) );
  CIVX2 U10 ( .A(c_out11), .Z(n3) );
  CIVX2 U11 ( .A(s2), .Z(n5) );
  CMXI2X1 U12 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_2841 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2842 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1421 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2842 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2841 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2843 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2844 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1422 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2844 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2843 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2845 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n4;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(n2) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U4 ( .A(b), .Z(n4) );
  CENX1 U5 ( .A(n4), .B(n2), .Z(sum) );
endmodule


module Add_half_2846 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVX1 U1 ( .A(b), .Z(n2) );
  CND2X1 U2 ( .A(n1), .B(b), .Z(n4) );
  CIVX1 U3 ( .A(a), .Z(n1) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CND2XL U5 ( .A(a), .B(n2), .Z(n3) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1423 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2846 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2845 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2847 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2848 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1424 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2848 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2847 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_356 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1424 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1423 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1422 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1421 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n2) );
  CMX2XL U4 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CMXI2X1 U5 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n3) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(c_out10), .Z(n5) );
  CIVX2 U10 ( .A(c_out11), .Z(n4) );
endmodule


module bit4_89 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_356 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_355 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_354 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_353 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVDX1 U3 ( .A(n8), .Z0(n1), .Z1(n2) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(c_out4) );
  CMX2XL U5 ( .A0(s43[0]), .A1(s44[0]), .S(n8), .Z(sum4[2]) );
  CND2XL U6 ( .A(c_out411), .B(n8), .Z(n4) );
  CMXI2X1 U7 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n5) );
  CIVX2 U8 ( .A(n5), .Z(n8) );
  CMX2X1 U9 ( .A0(s43[1]), .A1(s44[1]), .S(n2), .Z(sum4[3]) );
  CND2X1 U10 ( .A(c_out410), .B(n1), .Z(n3) );
  CMX2X1 U11 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U12 ( .A(s41[1]), .Z(n7) );
  CIVX2 U13 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
endmodule


module Add_half_2849 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2850 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1425 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2850 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2849 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2851 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2852 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1426 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2852 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2851 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2853 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2854 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1427 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2854 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2853 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2855 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2856 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1428 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2856 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2855 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_357 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1428 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1427 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1426 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1425 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_2857 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2858 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1429 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2858 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2857 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2859 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2860 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1430 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2860 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2859 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2861 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2862 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1431 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2862 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2861 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2863 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2864 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1432 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2864 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2863 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_358 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1432 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1431 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1430 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1429 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_2865 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2866 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1433 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2866 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2865 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2867 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2868 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1434 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2868 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2867 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2869 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2870 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1435 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2870 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2869 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2871 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2872 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1436 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2872 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2871 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_359 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1436 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1435 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1434 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1433 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n4), .S(n1), .Z(c_out2) );
  CMXI2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n4) );
  CIVX2 U8 ( .A(c_out11), .Z(n3) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_2873 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2874 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1437 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2874 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2873 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2875 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2876 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1438 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2876 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2875 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2877 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2878 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1439 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2878 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2877 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2879 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2880 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1440 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2880 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2879 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_360 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1440 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1439 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1438 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1437 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_90 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_360 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_359 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_358 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_357 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(c_in4), .Z(n2) );
  CMXI2X1 U4 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out4) );
  CIVDXL U5 ( .A(n3), .Z0(n10) );
  CIVX1 U6 ( .A(s41[0]), .Z(n7) );
  CMXI2X1 U7 ( .A0(c_out401), .A1(c_out400), .S(n2), .Z(n3) );
  CIVX1 U8 ( .A(s42[0]), .Z(n6) );
  CMXI2XL U9 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CMXI2XL U10 ( .A0(n12), .A1(n11), .S(n10), .Z(sum4[3]) );
  CMX2X1 U11 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(c_out410), .Z(n5) );
  CIVX2 U13 ( .A(c_out411), .Z(n4) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U15 ( .A(s43[0]), .Z(n9) );
  CIVX2 U16 ( .A(s44[0]), .Z(n8) );
  CIVX2 U17 ( .A(s43[1]), .Z(n12) );
  CIVX2 U18 ( .A(s44[1]), .Z(n11) );
endmodule


module Add_half_2881 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2882 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1441 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2882 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2881 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2883 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2884 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1442 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2884 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2883 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2885 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2886 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1443 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2886 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2885 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2887 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2888 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1444 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2888 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2887 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_361 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1444 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1443 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1442 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1441 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n7), .A1(n6), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n7) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
endmodule


module Add_half_2889 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2890 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1445 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2890 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2889 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2891 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2892 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1446 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2892 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2891 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2893 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2894 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1447 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2894 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2893 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2895 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2896 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1448 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2896 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2895 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_362 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1448 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1447 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1446 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1445 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
endmodule


module Add_half_2897 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2898 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1449 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2898 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2897 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2899 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2900 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1450 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2900 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2899 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2901 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2902 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1451 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2902 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2901 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2903 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2904 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1452 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2904 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2903 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_363 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1452 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1451 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1450 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1449 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_2905 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2906 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1453 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2906 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2905 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2907 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2908 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1454 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2908 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2907 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2909 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2910 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1455 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2910 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2909 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2911 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2912 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1456 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2912 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2911 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_364 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1456 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1455 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1454 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1453 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_91 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_364 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_363 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_362 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_361 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(n2), .Z(n1) );
  CMX2XL U4 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2XL U5 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U7 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX1 U8 ( .A(c_out411), .Z(n3) );
  CIVX1 U9 ( .A(c_out410), .Z(n4) );
  CMXI2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CMXI2X1 U11 ( .A0(n4), .A1(n3), .S(n1), .Z(c_out4) );
endmodule


module Add_half_2913 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2914 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1457 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2914 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2913 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2915 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2916 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1458 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2916 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2915 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2917 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2918 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1459 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2918 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2917 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2919 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2920 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1460 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2920 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2919 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_365 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1460 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1459 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1458 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1457 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2921 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2922 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1461 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2922 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2921 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2923 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2924 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1462 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2924 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2923 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2925 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2926 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1463 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2926 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2925 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2927 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2928 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1464 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2928 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2927 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_366 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1464 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1463 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1462 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1461 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2929 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2930 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1465 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2930 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2929 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2931 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2932 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1466 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2932 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2931 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2933 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2934 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1467 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2934 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2933 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2935 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2936 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1468 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2936 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2935 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_367 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1468 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1467 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1466 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1465 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U4 ( .A(c_out10), .Z(n3) );
  CIVX1 U5 ( .A(n1), .Z(n4) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2937 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2938 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1469 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2938 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2937 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2939 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2940 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1470 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2940 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2939 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2941 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2942 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1471 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2942 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2941 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2943 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2944 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1472 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2944 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2943 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_368 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1472 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1471 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1470 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1469 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_92 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_368 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_367 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_366 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_365 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(c_out411), .Z(n2) );
  CIVXL U4 ( .A(s43[1]), .Z(n12) );
  CMXI2XL U5 ( .A0(n12), .A1(n11), .S(n10), .Z(sum4[3]) );
  CMXI2XL U6 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n10) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n10), .Z(c_out4) );
  CIVX2 U11 ( .A(s41[0]), .Z(n5) );
  CIVX2 U12 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U14 ( .A(s41[1]), .Z(n7) );
  CIVX2 U15 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U16 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U17 ( .A(s43[0]), .Z(n9) );
  CIVX2 U18 ( .A(s44[0]), .Z(n8) );
  CIVX2 U19 ( .A(s44[1]), .Z(n11) );
endmodule


module bit8_23 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   n7, c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n5, n6;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_92 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_91 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_90 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_89 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X1 U3 ( .A0(s83[0]), .A1(s84[0]), .S(n6), .Z(sum8[4]) );
  CNIVX2 U4 ( .A(n6), .Z(n2) );
  CMX2X1 U5 ( .A0(c_out811), .A1(c_out810), .S(n3), .Z(c_out8) );
  CIVX1 U6 ( .A(n3), .Z(n1) );
  CMX2X2 U7 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2X1 U8 ( .A0(s83[3]), .A1(s84[3]), .S(n2), .Z(sum8[7]) );
  CNIVX3 U9 ( .A(n7), .Z(sum8[1]) );
  CMX2X2 U10 ( .A0(s81[0]), .A1(s82[0]), .S(c_in8), .Z(sum8[0]) );
  CIVX2 U11 ( .A(n5), .Z(n6) );
  CMX2XL U12 ( .A0(s83[1]), .A1(s84[1]), .S(n1), .Z(sum8[5]) );
  CMXI2X1 U13 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n3) );
  CMX2X2 U14 ( .A0(s83[2]), .A1(s84[2]), .S(n2), .Z(sum8[6]) );
  CMX2XL U15 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2XL U16 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(n7) );
  CMXI2X1 U17 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n5) );
endmodule


module Add_half_2945 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2946 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1473 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2946 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2945 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_2947 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2948 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1474 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2948 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2947 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2949 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2950 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1475 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2950 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2949 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_2951 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2952 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X2 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1476 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2952 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2951 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_369 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1476 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1475 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1474 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1473 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(n6), .Z(n1) );
  CIVXL U4 ( .A(n1), .Z(n2) );
  CMXI2XL U5 ( .A0(n8), .A1(n7), .S(n2), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(c_out10), .A1(c_out11), .S(n6), .Z(c_out2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CIVX2 U8 ( .A(n3), .Z(n6) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s3), .Z(n8) );
  CIVX2 U13 ( .A(s4), .Z(n7) );
endmodule


module Add_half_2953 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2954 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1477 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2954 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2953 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2955 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2956 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1478 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2956 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2955 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2957 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(a), .B(n2), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_2958 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1479 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2958 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2957 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2959 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2960 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1480 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2960 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2959 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_370 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1480 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1479 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1478 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1477 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2961 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2962 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1481 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2962 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2961 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2963 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2964 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1482 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2964 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2963 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2965 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2966 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1483 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2966 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2965 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_2967 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2968 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1484 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2968 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2967 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_371 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1484 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1483 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1482 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1481 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_2969 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2970 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1485 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2970 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2969 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2971 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2972 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1486 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2972 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2971 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2973 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2974 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1487 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_2974 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2973 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_2975 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2976 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1488 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2976 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2975 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_372 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1488 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1487 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1486 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1485 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_93 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_372 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_371 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_370 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_369 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n6), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n6), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(c_out410), .A1(c_out411), .S(n6), .Z(c_out4) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CIVX2 U8 ( .A(s41[0]), .Z(n3) );
  CIVX2 U9 ( .A(s42[0]), .Z(n2) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U11 ( .A(s41[1]), .Z(n5) );
  CIVX2 U12 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
endmodule


module Add_half_2977 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2978 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1489 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2978 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2977 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2979 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2980 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1490 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2980 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2979 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2981 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2982 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1491 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2982 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2981 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2983 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2984 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1492 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2984 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2983 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_373 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1492 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1491 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1490 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1489 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out11), .A1(c_out10), .S(n1), .Z(c_out2) );
  CIVXL U4 ( .A(n1), .Z(n2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_2985 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2986 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1493 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2986 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2985 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2987 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2988 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1494 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2988 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2987 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2989 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_2990 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1495 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2990 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2989 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_2991 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_2992 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1496 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_2992 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2991 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_374 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1496 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1495 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1494 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1493 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_2993 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_2994 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1497 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2994 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2993 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2995 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_2996 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1498 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2996 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2995 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2997 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_2998 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_full_1499 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_2998 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2997 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_2999 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3000 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_full_1500 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3000 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_2999 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_375 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1500 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1499 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1498 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1497 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U7 ( .A(s1), .Z(n5) );
  CIVX2 U8 ( .A(s2), .Z(n4) );
  CMXI2X1 U9 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U10 ( .A(s3), .Z(n7) );
  CIVX2 U11 ( .A(s4), .Z(n6) );
  CMXI2X1 U12 ( .A0(n7), .A1(n6), .S(n1), .Z(sum2[1]) );
endmodule


module Add_half_3001 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3002 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1501 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3002 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3001 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3003 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3004 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1502 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3004 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3003 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3005 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3006 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_full_1503 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3006 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3005 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3007 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3008 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1504 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3008 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3007 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_376 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1504 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1503 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1502 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1501 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_94 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_376 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_375 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_374 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_373 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U4 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX1 U5 ( .A(s43[1]), .Z(n8) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n6) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out4) );
  CIVX2 U11 ( .A(s43[0]), .Z(n5) );
  CIVX2 U12 ( .A(s44[0]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(n6), .Z(sum4[2]) );
  CIVX2 U14 ( .A(s44[1]), .Z(n7) );
  CMXI2X1 U15 ( .A0(n8), .A1(n7), .S(n6), .Z(sum4[3]) );
endmodule


module Add_half_3009 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3010 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1505 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3010 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3009 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3011 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3012 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1506 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3012 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3011 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3013 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3014 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1507 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3014 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3013 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3015 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3016 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1508 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3016 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3015 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_377 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1508 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1507 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1506 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1505 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3017 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3018 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1509 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3018 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3017 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3019 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3020 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1510 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3020 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3019 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3021 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3022 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1511 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3022 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3021 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3023 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3024 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1512 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3024 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3023 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_378 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1512 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1511 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1510 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1509 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3025 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3026 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1513 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3026 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3025 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3027 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3028 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1514 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3028 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3027 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3029 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3030 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1515 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3030 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3029 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3031 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3032 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1516 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3032 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3031 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_379 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1516 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1515 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1514 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1513 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3033 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3034 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1517 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3034 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3033 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3035 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3036 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1518 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3036 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3035 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3037 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3038 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1519 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3038 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3037 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3039 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3040 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1520 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3040 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3039 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_380 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1520 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1519 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1518 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1517 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_95 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_380 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_379 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_378 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_377 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_3041 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3042 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1521 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3042 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3041 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3043 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3044 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1522 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3044 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3043 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3045 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3046 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1523 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3046 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3045 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3047 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3048 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1524 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3048 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3047 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_381 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1524 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1523 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1522 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1521 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3049 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3050 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1525 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3050 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3049 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3051 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3052 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1526 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3052 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3051 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3053 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3054 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1527 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3054 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3053 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3055 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3056 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1528 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3056 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3055 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_382 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1528 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1527 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1526 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1525 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3057 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3058 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1529 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3058 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3057 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3059 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3060 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1530 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3060 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3059 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3061 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3062 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1531 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3062 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3061 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3063 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3064 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1532 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3064 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3063 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_383 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1532 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1531 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1530 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1529 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3065 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3066 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1533 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3066 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3065 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3067 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3068 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1534 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3068 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3067 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3069 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3070 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1535 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3070 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3069 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3071 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3072 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1536 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3072 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3071 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_384 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1536 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1535 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1534 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1533 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_96 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_384 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_383 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_382 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_381 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_24 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_96 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_95 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_94 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_93 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n3), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n3), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n3), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n3), .Z(sum8[0]) );
  CMX2X2 U3 ( .A0(s83[2]), .A1(s84[2]), .S(n1), .Z(sum8[6]) );
  CMX2X2 U4 ( .A0(s83[0]), .A1(s84[0]), .S(n1), .Z(sum8[4]) );
  CMX2X1 U5 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CMXI2X1 U6 ( .A0(c_out810), .A1(c_out811), .S(n1), .Z(n2) );
  CIVX2 U7 ( .A(n2), .Z(c_out8) );
  CMX2X2 U8 ( .A0(s83[3]), .A1(s84[3]), .S(n1), .Z(sum8[7]) );
  CMX2X2 U9 ( .A0(s83[1]), .A1(s84[1]), .S(n1), .Z(sum8[5]) );
  CIVX2 U14 ( .A(c_in8), .Z(n3) );
endmodule


module bit32_6 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   c1, c2, c3, n1, n2, n3, n4, n5;

  bit8_24 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8({a32[7], n3, a32[5:0]}), 
        .b8(b32[7:0]), .c_in8(c_in32) );
  bit8_23 A322 ( .sum8(sum32[15:8]), .c_out8(c2), .a8({a32[15:13], n5, 
        a32[11:9], n1}), .b8(b32[15:8]), .c_in8(c1) );
  bit8_22 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8(a32[23:16]), .b8(
        b32[23:16]), .c_in8(c2) );
  bit8_21 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8(a32[31:24]), .b8(
        b32[31:24]), .c_in8(c3) );
  CIVX4 U1 ( .A(n4), .Z(n5) );
  CIVX1 U2 ( .A(a32[6]), .Z(n2) );
  CNIVX4 U3 ( .A(a32[8]), .Z(n1) );
  CIVX4 U4 ( .A(n2), .Z(n3) );
  CIVX2 U5 ( .A(a32[12]), .Z(n4) );
endmodule


module Add_half_3073 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3074 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1537 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3074 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3073 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3075 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3076 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1538 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3076 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3075 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3077 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3078 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1539 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3078 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3077 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3079 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3080 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1540 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3080 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3079 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_385 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1540 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1539 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1538 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1537 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CIVX1 U5 ( .A(s4), .Z(n4) );
  CIVX2 U6 ( .A(s1), .Z(n3) );
  CIVX2 U7 ( .A(s2), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
endmodule


module Add_half_3081 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3082 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1541 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3082 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3081 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3083 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3084 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1542 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3084 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3083 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3085 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3086 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1543 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3086 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3085 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3087 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3088 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1544 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3088 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3087 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_386 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_1544 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1543 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1542 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1541 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(s3), .Z(n3) );
  CIVX2 U7 ( .A(s4), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(sum2[1]) );
endmodule


module Add_half_3089 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3090 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1545 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3090 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3089 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3091 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3092 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1546 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3092 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3091 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3093 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3094 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1547 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3094 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3093 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3095 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3096 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1548 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3096 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3095 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_387 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1548 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1547 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1546 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1545 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n6) );
  CMXI2X1 U4 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3097 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3098 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1549 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3098 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3097 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3099 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3100 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1550 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3100 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3099 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3101 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3102 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1551 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3102 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3101 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3103 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3104 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1552 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3104 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3103 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_388 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1552 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1551 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1550 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1549 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX1 U4 ( .A(n1), .Z(n4) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module bit4_97 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_388 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_387 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_386 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_385 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U7 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMX2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
endmodule


module Add_half_3105 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3106 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1553 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3106 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3105 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3107 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3108 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1554 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3108 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3107 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3109 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3110 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1555 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3110 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3109 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3111 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3112 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1556 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3112 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3111 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_389 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1;

  Add_full_1556 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1555 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1554 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1553 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3113 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3114 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1557 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3114 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3113 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3115 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3116 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1558 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3116 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3115 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3117 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3118 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1559 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3118 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3117 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3119 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3120 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1560 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3120 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3119 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_390 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1;

  Add_full_1560 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1559 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1558 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1557 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3121 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3122 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1561 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3122 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3121 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3123 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3124 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1562 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3124 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3123 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3125 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3126 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1563 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3126 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3125 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3127 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3128 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1564 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3128 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3127 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_391 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1564 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1563 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1562 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1561 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2X1 U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_3129 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3130 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1565 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3130 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3129 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3131 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3132 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1566 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3132 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3131 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3133 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3134 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1567 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3134 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3133 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3135 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3136 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1568 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3136 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3135 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_392 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1568 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1567 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1566 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1565 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n4) );
endmodule


module bit4_98 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_392 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_391 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_390 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_389 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMX2XL U4 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CIVX2 U6 ( .A(s41[0]), .Z(n3) );
  CIVX2 U7 ( .A(s42[0]), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U9 ( .A(s41[1]), .Z(n5) );
  CIVX2 U10 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(s43[0]), .Z(n7) );
  CIVX2 U13 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n1), .Z(sum4[2]) );
endmodule


module Add_half_3137 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3138 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1569 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3138 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3137 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3139 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3140 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1570 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3140 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3139 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3141 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3142 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1571 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3142 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3141 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3143 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3144 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1572 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3144 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3143 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_393 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1572 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1571 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1570 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1569 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U5 ( .A(s1), .Z(n3) );
  CMX2X1 U6 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CIVX2 U7 ( .A(s2), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
endmodule


module Add_half_3145 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3146 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1573 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3146 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3145 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3147 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3148 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1574 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3148 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3147 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3149 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3150 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1575 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3150 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3149 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3151 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3152 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1576 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3152 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3151 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_394 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1;

  Add_full_1576 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1575 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1574 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1573 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3153 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3154 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1577 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3154 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3153 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3155 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3156 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1578 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3156 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3155 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3157 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3158 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1579 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3158 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3157 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3159 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3160 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1580 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3160 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3159 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_395 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1580 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1579 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1578 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1577 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMX2X1 U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMXI2X1 U5 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n3) );
  CMX2XL U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMXI2X1 U7 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CIVX1 U8 ( .A(s2), .Z(n6) );
  CIVX1 U9 ( .A(s1), .Z(n7) );
  CIVX2 U10 ( .A(c_out10), .Z(n5) );
  CIVX2 U11 ( .A(c_out11), .Z(n4) );
  CMXI2X1 U12 ( .A0(n7), .A1(n6), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3161 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3162 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1581 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3162 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3161 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3163 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3164 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1582 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3164 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3163 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3165 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3166 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1583 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3166 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3165 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3167 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3168 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n1), .B(b), .Z(n4) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1584 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3168 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3167 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_396 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1584 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1583 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1582 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1581 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n3) );
  CMX2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMXI2X1 U6 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(c_out10), .Z(n5) );
  CIVX2 U10 ( .A(c_out11), .Z(n4) );
endmodule


module bit4_99 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_396 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_395 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_394 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_393 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(c_in4), .Z(n2) );
  CIVX2 U4 ( .A(n3), .Z(n1) );
  CMXI2X1 U5 ( .A0(c_out401), .A1(c_out400), .S(n2), .Z(n3) );
  CIVX1 U6 ( .A(s42[1]), .Z(n6) );
  CMX2XL U7 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U8 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U9 ( .A(c_out410), .Z(n5) );
  CIVX2 U10 ( .A(c_out411), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(n1), .Z(c_out4) );
  CIVX2 U12 ( .A(s41[1]), .Z(n7) );
  CMXI2X1 U13 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n9) );
  CIVX2 U15 ( .A(s44[0]), .Z(n8) );
  CMXI2X1 U16 ( .A0(n9), .A1(n8), .S(n1), .Z(sum4[2]) );
endmodule


module Add_half_3169 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3170 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1585 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3170 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3169 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3171 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3172 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1586 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3172 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3171 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3173 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3174 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1587 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3174 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3173 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3175 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3176 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1588 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3176 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3175 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_397 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1;

  Add_full_1588 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1587 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1586 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1585 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2X1 U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3177 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3178 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1589 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3178 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3177 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3179 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3180 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1590 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3180 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3179 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3181 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3182 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1591 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3182 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3181 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3183 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3184 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1592 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3184 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3183 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_398 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1;

  Add_full_1592 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1591 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1590 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1589 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3185 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3186 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1593 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3186 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3185 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3187 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3188 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1594 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3188 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3187 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3189 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n3;

  CENX1 U1 ( .A(n3), .B(n1), .Z(sum) );
  CNIVXL U2 ( .A(a), .Z(n1) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U4 ( .A(b), .Z(n3) );
endmodule


module Add_half_3190 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1595 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3190 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3189 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3191 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(n1), .Z(sum) );
endmodule


module Add_half_3192 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1596 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3192 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3191 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_399 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1596 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1595 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1594 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1593 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n2), .Z(n7) );
  CIVXL U4 ( .A(s1), .Z(n6) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U6 ( .A0(n3), .A1(n4), .S(n1), .Z(c_out2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMX2XL U8 ( .A0(s3), .A1(s4), .S(n7), .Z(sum2[1]) );
  CIVX1 U9 ( .A(s2), .Z(n5) );
  CIVX2 U10 ( .A(c_out10), .Z(n4) );
  CIVX2 U11 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U12 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3193 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3194 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1597 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3194 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3193 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3195 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3196 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1598 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3196 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3195 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3197 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3198 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1599 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3198 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3197 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3199 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3200 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n1), .B(b), .Z(n4) );
  CIVX1 U2 ( .A(a), .Z(n1) );
  CND2XL U3 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1600 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3200 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3199 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_400 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1600 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1599 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1598 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1597 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMXI2XL U5 ( .A0(n6), .A1(n5), .S(n1), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n4) );
  CIVX2 U8 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module bit4_100 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_400 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_399 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_398 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_397 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(s44[0]), .Z(n4) );
  CIVX2 U4 ( .A(n1), .Z(n6) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2X1 U6 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out4) );
  CMX2XL U7 ( .A0(s43[1]), .A1(s44[1]), .S(n6), .Z(sum4[3]) );
  CMX2X1 U8 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U9 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX1 U10 ( .A(c_out410), .Z(n3) );
  CIVX2 U11 ( .A(c_out411), .Z(n2) );
  CIVX2 U12 ( .A(s43[0]), .Z(n5) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(n6), .Z(sum4[2]) );
endmodule


module bit8_25 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   n31, c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n23, n24, n25, n26, n27, n28, n29, n30;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_100 A81 ( .sum4(s81), .c_out4(c_out800), .a4({a8[3:1], n24}), .b4(
        b8[3:0]), .c_in4(1'b0) );
  bit4_99 A82 ( .sum4(s82), .c_out4(c_out801), .a4({a8[3:1], n24}), .b4(
        b8[3:0]), .c_in4(1'b1) );
  bit4_98 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_97 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVX3 U3 ( .A(n20), .Z(n17) );
  CND2X4 U4 ( .A(n17), .B(s83[0]), .Z(n15) );
  CND2X2 U5 ( .A(c_out801), .B(n6), .Z(n10) );
  CIVX2 U6 ( .A(n1), .Z(sum8[1]) );
  CIVX4 U7 ( .A(n23), .Z(n24) );
  CND2X1 U8 ( .A(s84[3]), .B(n7), .Z(n14) );
  CMXI2X1 U9 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(n1) );
  CIVX1 U10 ( .A(n20), .Z(n2) );
  CND2X4 U11 ( .A(n11), .B(n12), .Z(sum8[5]) );
  CND2X2 U12 ( .A(s82[2]), .B(n3), .Z(n4) );
  CND2X1 U13 ( .A(s81[2]), .B(n8), .Z(n5) );
  CND2X4 U14 ( .A(n4), .B(n5), .Z(sum8[2]) );
  CIVX1 U15 ( .A(n8), .Z(n3) );
  CND2X4 U16 ( .A(n18), .B(n19), .Z(sum8[6]) );
  CNIVX1 U17 ( .A(c_in8), .Z(n6) );
  CIVX1 U18 ( .A(c_in8), .Z(n8) );
  CIVX1 U19 ( .A(s82[3]), .Z(n29) );
  CND2X1 U20 ( .A(s84[1]), .B(n20), .Z(n12) );
  CND2X2 U21 ( .A(s84[0]), .B(n20), .Z(n16) );
  CND2X1 U22 ( .A(s84[2]), .B(n20), .Z(n19) );
  CIVXL U23 ( .A(n2), .Z(n7) );
  CND2X1 U24 ( .A(c_out800), .B(n8), .Z(n9) );
  CND2X2 U25 ( .A(n9), .B(n10), .Z(n20) );
  CIVX1 U26 ( .A(s81[3]), .Z(n30) );
  CMXI2XL U27 ( .A0(n26), .A1(n25), .S(n7), .Z(c_out8) );
  CND2X1 U28 ( .A(s83[1]), .B(n2), .Z(n11) );
  CND2X2 U29 ( .A(n13), .B(n14), .Z(sum8[7]) );
  CND2X1 U30 ( .A(s83[3]), .B(n2), .Z(n13) );
  CMXI2X1 U31 ( .A0(n30), .A1(n29), .S(n3), .Z(n31) );
  CIVX2 U32 ( .A(n31), .Z(n21) );
  CND2X1 U33 ( .A(s83[2]), .B(n2), .Z(n18) );
  CND2X4 U34 ( .A(n15), .B(n16), .Z(sum8[4]) );
  CIVX4 U35 ( .A(n21), .Z(sum8[3]) );
  CIVX1 U36 ( .A(s81[0]), .Z(n28) );
  CIVX2 U37 ( .A(a8[0]), .Z(n23) );
  CMXI2X1 U38 ( .A0(n28), .A1(n27), .S(c_in8), .Z(sum8[0]) );
  CIVX2 U39 ( .A(c_out810), .Z(n26) );
  CIVX2 U40 ( .A(c_out811), .Z(n25) );
  CIVX2 U41 ( .A(s82[0]), .Z(n27) );
endmodule


module Add_half_3201 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3202 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1601 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3202 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3201 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3203 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3204 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1602 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3204 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3203 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3205 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOX2 U1 ( .A(b), .B(n1), .Z(sum) );
  CNIVX1 U2 ( .A(a), .Z(n1) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3206 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1603 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3206 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3205 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3207 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3208 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1604 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3208 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3207 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_401 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1604 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1603 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1602 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1601 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n4), .A1(n3), .S(n1), .Z(c_out2) );
  CMXI2XL U4 ( .A0(n6), .A1(n5), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out10), .Z(n4) );
  CIVX2 U9 ( .A(c_out11), .Z(n3) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module Add_half_3209 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3210 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1605 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3210 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3209 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3211 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3212 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1606 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3212 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3211 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3213 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3214 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1607 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3214 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3213 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3215 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3216 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1608 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3216 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3215 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_402 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_1608 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1607 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1606 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1605 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U5 ( .A(c_out10), .Z(n3) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
endmodule


module Add_half_3217 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3218 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1609 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3218 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3217 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3219 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3220 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1610 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3220 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3219 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3221 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3222 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1611 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3222 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3221 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3223 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3224 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1612 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3224 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3223 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_403 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1612 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1611 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1610 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1609 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CIVX2 U4 ( .A(n1), .Z(n6) );
  CIVX1 U5 ( .A(s2), .Z(n4) );
  CIVX1 U6 ( .A(s1), .Z(n5) );
  CIVX1 U7 ( .A(c_out10), .Z(n3) );
  CIVX1 U8 ( .A(c_out11), .Z(n2) );
  CMXI2XL U9 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
  CMXI2X1 U10 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s3), .Z(n8) );
  CIVX2 U13 ( .A(s4), .Z(n7) );
endmodule


module Add_half_3225 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3226 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1613 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3226 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3225 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3227 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3228 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1614 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3228 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3227 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3229 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3230 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1615 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3230 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3229 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3231 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3232 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(b), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U3 ( .A(b), .Z(n1) );
  CIVX1 U4 ( .A(a), .Z(n2) );
  CND2X1 U5 ( .A(n1), .B(a), .Z(n4) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1616 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3232 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3231 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_404 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1616 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1615 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1614 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1613 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(n2), .Z(n5) );
  CMXI2X1 U4 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CIVX20 U6 ( .A(c_in2), .Z(n1) );
  CIVX1 U7 ( .A(c_out10), .Z(n4) );
  CIVX1 U8 ( .A(c_out11), .Z(n3) );
  CMX2XL U9 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U10 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module bit4_101 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_404 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_403 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_402 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_401 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CNIVX2 U3 ( .A(n8), .Z(n4) );
  CND2XL U4 ( .A(c_out410), .B(n1), .Z(n2) );
  CND2XL U5 ( .A(c_out411), .B(n8), .Z(n3) );
  CND2X1 U6 ( .A(n2), .B(n3), .Z(c_out4) );
  CIVXL U7 ( .A(n8), .Z(n1) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n5) );
  CMX2X1 U9 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMXI2X1 U10 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX1 U11 ( .A(s44[0]), .Z(n6) );
  CMX2X1 U12 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U13 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U14 ( .A(n5), .Z(n8) );
  CIVX2 U15 ( .A(s43[0]), .Z(n7) );
endmodule


module Add_half_3233 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3234 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1617 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3234 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3233 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3235 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3236 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1618 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3236 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3235 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3237 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3238 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1619 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3238 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3237 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3239 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3240 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n3), .B(n4), .Z(sum) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n1), .B(b), .Z(n4) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1620 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3240 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3239 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_405 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1620 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1619 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1618 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1617 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CIVX2 U4 ( .A(c_in2), .Z(n2) );
  CMXI2XL U5 ( .A0(n8), .A1(n7), .S(n1), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_out10), .Z(n4) );
  CIVX2 U7 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U8 ( .A0(n4), .A1(n3), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n6) );
  CIVX2 U10 ( .A(s2), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s3), .Z(n8) );
  CIVX2 U13 ( .A(s4), .Z(n7) );
endmodule


module Add_half_3241 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(a), .B(n2), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3242 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1621 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3242 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3241 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3243 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3244 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1622 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3244 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3243 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3245 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3246 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1623 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3246 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3245 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3247 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3248 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1624 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3248 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3247 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_406 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1624 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1623 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1622 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1621 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_3249 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3250 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1625 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3250 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3249 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3251 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3252 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1626 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3252 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3251 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3253 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3254 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1627 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3254 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3253 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3255 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3256 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1628 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3256 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3255 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_407 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1628 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1627 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1626 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1625 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n2), .Z(n7) );
  CIVX2 U4 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U5 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CIVX2 U6 ( .A(c_out11), .Z(n3) );
  CIVX1 U7 ( .A(s1), .Z(n6) );
  CIVX2 U8 ( .A(c_out10), .Z(n4) );
  CMX2XL U9 ( .A0(s3), .A1(s4), .S(n7), .Z(sum2[1]) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(n7), .Z(c_out2) );
  CIVX2 U11 ( .A(s2), .Z(n5) );
  CMXI2X1 U12 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3257 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3258 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1629 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3258 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3257 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3259 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3260 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1630 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3260 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3259 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3261 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3262 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1631 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3262 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3261 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3263 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3264 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1632 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3264 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3263 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_408 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1632 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1631 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1630 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1629 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n4) );
  CMXI2X1 U4 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX1 U5 ( .A(c_out11), .Z(n2) );
  CIVX1 U6 ( .A(c_out10), .Z(n3) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module bit4_102 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_408 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_407 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_406 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_405 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(c_out410), .A1(c_out411), .S(n4), .Z(c_out4) );
  CIVX2 U4 ( .A(n1), .Z(n4) );
  CMX2XL U5 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U7 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U9 ( .A(s41[1]), .Z(n3) );
  CIVX2 U10 ( .A(s42[1]), .Z(n2) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(c_in4), .Z(sum4[1]) );
endmodule


module Add_half_3265 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3266 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1633 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3266 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3265 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3267 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3268 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1634 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3268 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3267 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3269 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3270 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1635 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3270 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3269 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_3271 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3272 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2XL U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1636 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3272 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3271 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_409 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1636 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1635 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1634 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1633 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s2), .Z(n4) );
  CIVX1 U4 ( .A(s1), .Z(n5) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n6) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_3273 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3274 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1637 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3274 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3273 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3275 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3276 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1638 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3276 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3275 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3277 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3278 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1639 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3278 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3277 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3279 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CENXL U2 ( .A(a), .B(n2), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3280 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CIVX1 U1 ( .A(b), .Z(n2) );
  CENX1 U2 ( .A(a), .B(n2), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1640 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3280 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3279 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_410 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1640 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1639 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1638 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1637 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(n1), .Z(n4) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_3281 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3282 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(n1), .B(b), .Z(n4) );
  CIVXL U2 ( .A(a), .Z(n1) );
  CND2XL U3 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1641 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3282 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3281 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3283 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3284 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U2 ( .A(a), .B(n2), .Z(n3) );
  CIVXL U3 ( .A(a), .Z(n1) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1642 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3284 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3283 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3285 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENX1 U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3286 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(b), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n1), .B(a), .Z(n4) );
  CND2X2 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U4 ( .A(b), .Z(n1) );
  CIVX1 U5 ( .A(a), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1643 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3286 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3285 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3287 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3288 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n3), .B(n4), .Z(sum) );
  CND2X1 U2 ( .A(b), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n1), .B(a), .Z(n4) );
  CIVXL U4 ( .A(b), .Z(n1) );
  CIVX1 U5 ( .A(a), .Z(n2) );
  CAN2XL U6 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1644 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3288 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3287 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_411 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1644 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1643 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1642 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1641 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n2) );
  CIVX2 U4 ( .A(c_out11), .Z(n4) );
  CIVX1 U5 ( .A(c_out10), .Z(n5) );
  CMX2XL U6 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CMXI2X1 U7 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CMXI2X1 U8 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n3) );
  CMXI2XL U9 ( .A0(n7), .A1(n6), .S(n1), .Z(sum2[1]) );
  CMX2X1 U10 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n7) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
endmodule


module Add_half_3289 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3290 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(n1), .B(b), .Z(n4) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1645 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3290 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3289 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3291 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3292 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U2 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U3 ( .A(a), .Z(n1) );
  CND2X1 U4 ( .A(a), .B(n2), .Z(n3) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1646 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3292 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3291 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3293 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3294 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CIVX1 U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1647 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3294 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3293 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3295 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3296 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2, n3, n4, n5;

  CND2X1 U1 ( .A(n4), .B(n5), .Z(sum) );
  CND2X1 U2 ( .A(n2), .B(b), .Z(n5) );
  CIVDXL U3 ( .A(b), .Z0(n3) );
  CND2X1 U4 ( .A(a), .B(n3), .Z(n4) );
  CIVX1 U5 ( .A(a), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1648 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3296 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3295 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_412 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1648 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1647 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1646 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1645 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(c_out11), .Z(n3) );
  CIVX1 U4 ( .A(c_out10), .Z(n4) );
  CMX2XL U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U6 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module bit4_103 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_412 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_411 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_410 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_409 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X2 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX1 U4 ( .A(c_out410), .Z(n4) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CIVX1 U6 ( .A(c_out411), .Z(n3) );
  CMX2X1 U7 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CMXI2X1 U8 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out4) );
  CMX2XL U9 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U10 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U11 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
endmodule


module Add_half_3297 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3298 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1649 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3298 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3297 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3299 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3300 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1650 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3300 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3299 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3301 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3302 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1651 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3302 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3301 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3303 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3304 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1652 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3304 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3303 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_413 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1652 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1651 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1650 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1649 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_3305 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3306 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_full_1653 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3306 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3305 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3307 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(a), .B(n2), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3308 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1654 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3308 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3307 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3309 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3310 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1655 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3310 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3309 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3311 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3312 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1656 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3312 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3311 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_414 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1656 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1655 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1654 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1653 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n4) );
  CIVX2 U7 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n1), .Z(c_out2) );
endmodule


module Add_half_3313 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3314 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1657 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3314 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3313 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3315 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(a), .B(n2), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3316 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U2 ( .A(n3), .B(n4), .Z(sum) );
  CND2XL U3 ( .A(a), .B(n2), .Z(n3) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1658 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3316 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3315 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3317 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3318 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1659 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3318 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3317 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3319 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3320 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X2 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1660 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3320 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3319 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_415 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1660 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1659 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1658 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1657 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n3) );
  CMX2XL U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMXI2X1 U6 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CIVX1 U7 ( .A(s2), .Z(n6) );
  CIVX1 U8 ( .A(c_out10), .Z(n5) );
  CMX2XL U9 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_out11), .Z(n4) );
  CIVX2 U11 ( .A(s1), .Z(n7) );
  CMXI2X1 U12 ( .A0(n7), .A1(n6), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3321 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3322 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1661 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3322 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3321 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3323 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3324 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1662 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3324 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3323 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3325 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3326 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1663 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3326 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3325 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3327 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3328 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVX1 U1 ( .A(a), .Z(n1) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U4 ( .A(n4), .B(n3), .Z(sum) );
  CIVX1 U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1664 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3328 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3327 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_416 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1664 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1663 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1662 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1661 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out11), .Z(n3) );
  CIVX2 U4 ( .A(c_out10), .Z(n4) );
  CMX2XL U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U6 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module bit4_104 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_416 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_415 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_414 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_413 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n10), .A1(n9), .S(n1), .Z(sum4[3]) );
  CMX2X2 U4 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CIVX1 U6 ( .A(c_out411), .Z(n3) );
  CIVX1 U7 ( .A(c_out410), .Z(n4) );
  CIVX1 U8 ( .A(s43[0]), .Z(n8) );
  CIVX1 U9 ( .A(s44[0]), .Z(n7) );
  CMXI2X1 U10 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out4) );
  CMX2X1 U11 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX1 U12 ( .A(s44[1]), .Z(n9) );
  CIVX1 U13 ( .A(s43[1]), .Z(n10) );
  CIVX2 U14 ( .A(s41[1]), .Z(n6) );
  CIVX2 U15 ( .A(s42[1]), .Z(n5) );
  CMXI2X1 U16 ( .A0(n6), .A1(n5), .S(c_in4), .Z(sum4[1]) );
  CMXI2X1 U17 ( .A0(n8), .A1(n7), .S(n1), .Z(sum4[2]) );
endmodule


module bit8_26 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, net76382, net89774, net89773,
         net90251, net110968, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_104 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_103 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_102 A83 ( .sum4(s83), .c_out4(c_out810), .a4({a8[7], n14, n16, a8[4]}), 
        .b4({b8[7:6], n12, n20}), .c_in4(1'b0) );
  bit4_101 A84 ( .sum4(s84), .c_out4(c_out811), .a4({a8[7], n14, n5, a8[4]}), 
        .b4({b8[7:6], n1, n20}), .c_in4(1'b1) );
  CIVX1 U3 ( .A(s84[2]), .Z(n26) );
  CNIVX4 U4 ( .A(b8[5]), .Z(n1) );
  CND2X1 U5 ( .A(net89774), .B(net89773), .Z(n2) );
  CIVX2 U6 ( .A(n2), .Z(n11) );
  CND2X1 U7 ( .A(net89773), .B(net89774), .Z(n6) );
  CIVX2 U8 ( .A(a8[5]), .Z(n15) );
  CNIVX4 U9 ( .A(b8[4]), .Z(n20) );
  CIVX3 U10 ( .A(n15), .Z(n5) );
  CIVX2 U11 ( .A(net76382), .Z(net90251) );
  CND2IX1 U12 ( .B(n11), .A(c_out811), .Z(n9) );
  CMXI2X1 U13 ( .A0(n3), .A1(n4), .S(c_in8), .Z(sum8[0]) );
  CIVX2 U14 ( .A(s82[0]), .Z(n4) );
  CIVX2 U15 ( .A(s81[0]), .Z(n3) );
  CIVX1 U16 ( .A(c_in8), .Z(net76382) );
  CND2IX1 U17 ( .B(c_in8), .A(c_out800), .Z(net89773) );
  CND2X1 U18 ( .A(c_in8), .B(c_out801), .Z(net89774) );
  CIVXL U19 ( .A(n11), .Z(n19) );
  CIVX3 U20 ( .A(n15), .Z(n16) );
  CMXI2X1 U21 ( .A0(n21), .A1(n22), .S(n6), .Z(sum8[4]) );
  CND2X2 U22 ( .A(s81[2]), .B(net110968), .Z(n7) );
  CND2X1 U23 ( .A(s82[2]), .B(net90251), .Z(n8) );
  CND2X2 U24 ( .A(n7), .B(n8), .Z(sum8[2]) );
  CIVX2 U25 ( .A(net90251), .Z(net110968) );
  CND2X1 U26 ( .A(c_out810), .B(n11), .Z(n10) );
  CND2X2 U27 ( .A(n9), .B(n10), .Z(c_out8) );
  CMXI2X1 U28 ( .A0(n24), .A1(n23), .S(n11), .Z(sum8[5]) );
  CND2X2 U29 ( .A(n17), .B(n18), .Z(sum8[3]) );
  CMX2X2 U30 ( .A0(s82[1]), .A1(s81[1]), .S(net76382), .Z(sum8[1]) );
  CMX2X2 U31 ( .A0(s83[3]), .A1(s84[3]), .S(n19), .Z(sum8[7]) );
  CMXI2X1 U32 ( .A0(n26), .A1(n25), .S(n11), .Z(sum8[6]) );
  CNIVX4 U33 ( .A(b8[5]), .Z(n12) );
  CIVX1 U34 ( .A(s83[2]), .Z(n25) );
  CIVX2 U35 ( .A(a8[6]), .Z(n13) );
  CIVX4 U36 ( .A(n13), .Z(n14) );
  CND2XL U37 ( .A(s81[3]), .B(net76382), .Z(n17) );
  CND2XL U38 ( .A(s82[3]), .B(net90251), .Z(n18) );
  CIVX2 U39 ( .A(s84[0]), .Z(n22) );
  CIVX2 U40 ( .A(s83[0]), .Z(n21) );
  CIVX2 U41 ( .A(s84[1]), .Z(n24) );
  CIVX2 U42 ( .A(s83[1]), .Z(n23) );
endmodule


module Add_half_3329 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3330 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1665 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3330 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3329 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3331 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3332 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1666 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3332 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3331 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3333 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n3;

  CENX1 U1 ( .A(n3), .B(n1), .Z(sum) );
  CNIVXL U2 ( .A(a), .Z(n1) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U4 ( .A(b), .Z(n3) );
endmodule


module Add_half_3334 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1667 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3334 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3333 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3335 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3336 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1668 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3336 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3335 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_417 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1668 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1667 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1666 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1665 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_3337 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3338 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1669 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3338 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3337 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3339 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3340 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1670 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3340 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3339 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3341 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3342 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1671 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3342 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3341 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3343 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3344 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1672 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3344 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3343 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_418 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1672 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1671 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1670 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1669 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CIVX2 U4 ( .A(c_in2), .Z(n2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3345 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3346 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1673 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3346 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3345 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3347 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3348 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1674 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3348 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3347 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3349 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3350 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1675 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3350 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3349 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_3351 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3352 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1676 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3352 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3351 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_419 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n2, n3, n4, n5,
         n6, n7, n8, n9;

  Add_full_1676 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1675 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1674 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1673 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CIVDXL U4 ( .A(n2), .Z0(n7) );
  CIVX1 U5 ( .A(c_out11), .Z(n3) );
  CMXI2XL U6 ( .A0(n9), .A1(n8), .S(n7), .Z(sum2[1]) );
  CIVX1 U7 ( .A(c_out10), .Z(n4) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX2 U9 ( .A(s1), .Z(n6) );
  CIVX2 U10 ( .A(s2), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s3), .Z(n9) );
  CIVX2 U13 ( .A(s4), .Z(n8) );
endmodule


module Add_half_3353 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3354 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1677 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3354 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3353 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3355 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3356 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1678 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3356 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3355 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3357 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3358 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVX1 U1 ( .A(a), .Z(n2) );
  CND2X1 U2 ( .A(n3), .B(n4), .Z(sum) );
  CND2XL U3 ( .A(n1), .B(a), .Z(n4) );
  CND2XL U4 ( .A(b), .B(n2), .Z(n3) );
  CIVXL U5 ( .A(b), .Z(n1) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1679 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3358 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3357 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_3359 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3360 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1680 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3360 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3359 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_420 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n2, n3, n4, n5;

  Add_full_1680 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1679 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1678 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1677 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CIVDXL U4 ( .A(n2), .Z0(n5) );
  CIVX1 U5 ( .A(c_out11), .Z(n3) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out10), .Z(n4) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module bit4_105 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_420 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_419 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_418 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_417 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CNIVXL U3 ( .A(n2), .Z(n1) );
  CIVX2 U4 ( .A(c_out411), .Z(n5) );
  CIVX2 U5 ( .A(c_out410), .Z(n4) );
  CMXI2X1 U6 ( .A0(n8), .A1(n7), .S(n1), .Z(sum4[3]) );
  CANR2X1 U7 ( .A(c_out400), .B(n3), .C(c_out401), .D(c_in4), .Z(n2) );
  CANR2X1 U8 ( .A(c_out400), .B(n3), .C(c_in4), .D(c_out401), .Z(n6) );
  CMX2X1 U9 ( .A0(s44[0]), .A1(s43[0]), .S(n2), .Z(sum4[2]) );
  CMX2X1 U10 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U11 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(c_in4), .Z(n3) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(n6), .Z(c_out4) );
  CIVX2 U14 ( .A(s44[1]), .Z(n8) );
  CIVX2 U15 ( .A(s43[1]), .Z(n7) );
endmodule


module Add_half_3361 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3362 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1681 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3362 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3361 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3363 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3364 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1682 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3364 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3363 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3365 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3366 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1683 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3366 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3365 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3367 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3368 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1684 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3368 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3367 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_421 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1684 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1683 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1682 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1681 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_3369 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3370 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1685 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3370 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3369 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3371 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3372 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1686 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3372 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3371 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3373 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3374 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1687 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3374 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3373 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_3375 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3376 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1688 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3376 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3375 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_422 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1688 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1687 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1686 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1685 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U4 ( .A(s2), .Z(n4) );
  CIVX1 U5 ( .A(s1), .Z(n5) );
  CMXI2XL U6 ( .A0(n7), .A1(n6), .S(n1), .Z(sum2[1]) );
  CIVX2 U7 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n7) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
endmodule


module Add_half_3377 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CENX1 U4 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3378 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENX2 U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_full_1689 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3378 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3377 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_3379 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3380 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_full_1690 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3380 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3379 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_3381 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3382 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(b), .B(n2), .Z(n3) );
  CIVX2 U2 ( .A(a), .Z(n2) );
  CND2XL U3 ( .A(n1), .B(a), .Z(n4) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n1) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1691 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3382 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3381 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_3383 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3384 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(a), .Z(n1) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CENX1 U3 ( .A(b), .B(n1), .Z(sum) );
endmodule


module Add_full_1692 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3384 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3383 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_423 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1692 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1691 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1690 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1689 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_out10), .Z(n4) );
  CIVX2 U7 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX2 U9 ( .A(s1), .Z(n6) );
  CIVX2 U10 ( .A(s2), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3385 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3386 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_full_1693 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3386 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3385 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3387 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3388 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1694 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3388 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3387 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3389 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3390 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U2 ( .A(a), .Z(n2) );
  CND2XL U3 ( .A(b), .B(n2), .Z(n3) );
  CND2X1 U4 ( .A(n1), .B(a), .Z(n4) );
  CIVXL U5 ( .A(b), .Z(n1) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1695 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3390 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3389 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_3391 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3392 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1696 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3392 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3391 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_424 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1696 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1695 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1694 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1693 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2X1 U3 ( .A(c_out00), .B(n5), .Z(n3) );
  CND2X1 U4 ( .A(n2), .B(n3), .Z(n4) );
  CMX2X1 U5 ( .A0(s4), .A1(s3), .S(n1), .Z(sum2[1]) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n5), .Z(n1) );
  CMX2XL U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CND2X1 U8 ( .A(c_out01), .B(c_in2), .Z(n2) );
  CIVX2 U9 ( .A(c_in2), .Z(n5) );
  CIVX2 U10 ( .A(c_out10), .Z(n7) );
  CIVX2 U11 ( .A(c_out11), .Z(n6) );
  CMXI2X1 U12 ( .A0(n7), .A1(n6), .S(n4), .Z(c_out2) );
endmodule


module bit4_106 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_424 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_423 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_422 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_421 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2XL U3 ( .A(n3), .B(c_out400), .C(c_in4), .D(c_out401), .Z(n1) );
  CANR2X1 U4 ( .A(n3), .B(c_out400), .C(c_in4), .D(c_out401), .Z(n2) );
  CANR2X1 U5 ( .A(n3), .B(c_out400), .C(c_in4), .D(c_out401), .Z(n4) );
  CMX2X1 U6 ( .A0(s44[0]), .A1(s43[0]), .S(n2), .Z(sum4[2]) );
  CMX2X1 U7 ( .A0(c_out411), .A1(c_out410), .S(n4), .Z(c_out4) );
  CMX2XL U8 ( .A0(s44[1]), .A1(s43[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U9 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U10 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U11 ( .A(c_in4), .Z(n3) );
endmodule


module Add_half_3393 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3394 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1697 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3394 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3393 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3395 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3396 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1698 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3396 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3395 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3397 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3398 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1699 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3398 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3397 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_3399 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3400 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1700 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3400 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3399 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_425 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1700 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1699 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1698 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1697 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2X1 U3 ( .A(n5), .B(c_out11), .Z(n3) );
  CND2X2 U4 ( .A(c_out10), .B(n1), .Z(n2) );
  CND2X2 U5 ( .A(n2), .B(n3), .Z(c_out2) );
  CIVX2 U6 ( .A(n5), .Z(n1) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n4) );
  CMXI2XL U8 ( .A0(n7), .A1(n6), .S(n5), .Z(sum2[1]) );
  CIVX1 U9 ( .A(n4), .Z(n5) );
  CIVX1 U10 ( .A(s4), .Z(n6) );
  CIVX1 U11 ( .A(s3), .Z(n7) );
  CMX2X1 U12 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3401 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3402 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1701 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3402 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3401 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3403 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3404 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2, n3, n4, n5;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CND2XL U2 ( .A(a), .B(n3), .Z(n4) );
  CND2XL U3 ( .A(n2), .B(b), .Z(n5) );
  CND2X1 U4 ( .A(n4), .B(n5), .Z(sum) );
  CIVXL U5 ( .A(a), .Z(n2) );
  CIVXL U6 ( .A(b), .Z(n3) );
endmodule


module Add_full_1702 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3404 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3403 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3405 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3406 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CIVXL U1 ( .A(a), .Z(n1) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n1), .B(b), .Z(n4) );
  CND2X1 U4 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1703 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3406 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3405 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CND2X1 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_3407 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3408 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1704 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3408 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3407 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_426 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1704 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1703 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1702 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1701 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2X2 U3 ( .A(c_out10), .B(n1), .Z(n2) );
  CND2X1 U4 ( .A(n7), .B(c_out11), .Z(n3) );
  CND2X2 U5 ( .A(n2), .B(n3), .Z(c_out2) );
  CIVX2 U6 ( .A(n7), .Z(n1) );
  CIVX1 U7 ( .A(s2), .Z(n5) );
  CIVX1 U8 ( .A(s1), .Z(n6) );
  CIVX1 U9 ( .A(n4), .Z(n7) );
  CMX2XL U10 ( .A0(s3), .A1(s4), .S(n7), .Z(sum2[1]) );
  CMXI2X1 U11 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n4) );
  CMXI2X1 U12 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3409 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3410 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88196;
  assign c_out = net88196;

  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(net88196) );
endmodule


module Add_full_1705 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3410 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3409 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n1), .B(n2), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_3411 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3412 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1706 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3412 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3411 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3413 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3414 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1707 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3414 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3413 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3415 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net85686, net106258, net106259, n1, n2;
  assign c_out = net85686;

  CNR2X2 U1 ( .A(n1), .B(n2), .Z(net85686) );
  CIVX2 U2 ( .A(a), .Z(n1) );
  CIVX2 U3 ( .A(b), .Z(n2) );
  CIVXL U4 ( .A(a), .Z(net106258) );
  CEOX2 U5 ( .A(b), .B(net106259), .Z(sum) );
  CIVX1 U6 ( .A(net106258), .Z(net106259) );
endmodule


module Add_half_3416 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88011, n1, n2, n3, n4;
  assign c_out = net88011;

  CIVX2 U1 ( .A(a), .Z(n1) );
  CND2X2 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X2 U3 ( .A(n4), .B(n3), .Z(sum) );
  CAN2XL U4 ( .A(a), .B(b), .Z(net88011) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CND2X1 U6 ( .A(a), .B(n2), .Z(n3) );
endmodule


module Add_full_1708 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3416 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3415 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n1), .B(n2), .Z(c_out) );
  CIVXL U2 ( .A(w2), .Z(n2) );
  CIVX2 U3 ( .A(w3), .Z(n1) );
endmodule


module bit2_427 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, net76754,
         net76755, net113041, net113040, n1, n2, n3, n4, n5, n6, n7;

  Add_full_1708 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1707 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1706 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1705 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(c_out00), .Z(n1) );
  CIVXL U4 ( .A(n1), .Z(n2) );
  CMX2XL U5 ( .A0(c_out01), .A1(n2), .S(n5), .Z(n3) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n5), .Z(n4) );
  CMXI2X1 U7 ( .A0(net113040), .A1(net113041), .S(n4), .Z(c_out2) );
  CIVX2 U8 ( .A(c_in2), .Z(n5) );
  CMXI2X1 U9 ( .A0(net76754), .A1(net76755), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U10 ( .A(c_out10), .Z(net113041) );
  CIVX2 U11 ( .A(c_out11), .Z(net113040) );
  CIVX1 U12 ( .A(s2), .Z(net76755) );
  CMXI2XL U13 ( .A0(n7), .A1(n6), .S(n3), .Z(sum2[1]) );
  CIVX2 U14 ( .A(s1), .Z(net76754) );
  CIVX2 U15 ( .A(s3), .Z(n7) );
  CIVX2 U16 ( .A(s4), .Z(n6) );
endmodule


module Add_half_3417 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(n2) );
  CEOXL U3 ( .A(b), .B(n2), .Z(sum) );
  CAN2X1 U4 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3418 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88198;
  assign c_out = net88198;

  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(net88198) );
endmodule


module Add_full_1709 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3418 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3417 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w2), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n1) );
endmodule


module Add_half_3419 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3420 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4, n5;

  CIVXL U1 ( .A(n2), .Z(n1) );
  CIVX2 U2 ( .A(a), .Z(n2) );
  CND2X2 U3 ( .A(n5), .B(n4), .Z(sum) );
  CND2X1 U4 ( .A(n2), .B(b), .Z(n5) );
  CND2X1 U5 ( .A(a), .B(n3), .Z(n4) );
  CIVX1 U6 ( .A(b), .Z(n3) );
  CAN2XL U7 ( .A(n1), .B(b), .Z(c_out) );
endmodule


module Add_full_1710 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3420 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3419 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3421 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n3;

  CNIVX1 U1 ( .A(a), .Z(n1) );
  CENX1 U2 ( .A(n3), .B(n1), .Z(sum) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U4 ( .A(b), .Z(n3) );
endmodule


module Add_half_3422 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1711 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3422 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3421 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3423 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENXL U1 ( .A(b), .B(a), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(sum) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3424 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1712 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3424 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3423 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_428 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, net85280,
         net108940, net108939, n1, n2, n3;

  Add_full_1712 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1711 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1710 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1709 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(net85280) );
  CMXI2XL U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CMXI2X1 U5 ( .A0(n1), .A1(n2), .S(net85280), .Z(c_out2) );
  CIVX1 U6 ( .A(c_out10), .Z(n2) );
  CIVX2 U7 ( .A(c_out11), .Z(n1) );
  CMXI2X1 U8 ( .A0(net108939), .A1(net108940), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(s1), .Z(net108939) );
  CIVX2 U10 ( .A(s2), .Z(net108940) );
  CMX2X1 U11 ( .A0(s4), .A1(s3), .S(n3), .Z(sum2[1]) );
endmodule


module bit4_107 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, net106317, net107963,
         net76801, net76800, net90809, net87659, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_428 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_427 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_426 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_425 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CND2IX1 U3 ( .B(c_in4), .A(c_out400), .Z(n1) );
  CND2X1 U4 ( .A(c_out401), .B(c_in4), .Z(net90809) );
  CND2X2 U5 ( .A(net90809), .B(n1), .Z(net87659) );
  CMXI2X1 U6 ( .A0(net76800), .A1(net76801), .S(net87659), .Z(c_out4) );
  CND2X1 U7 ( .A(n1), .B(net90809), .Z(net107963) );
  CMX2X1 U8 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U9 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U10 ( .A(c_out411), .Z(net76801) );
  CIVX2 U11 ( .A(c_out410), .Z(net76800) );
  CIVX1 U12 ( .A(net107963), .Z(net106317) );
  CND2X1 U13 ( .A(s43[0]), .B(net106317), .Z(n2) );
  CND2XL U14 ( .A(net107963), .B(s44[0]), .Z(n3) );
  CND2X1 U15 ( .A(n2), .B(n3), .Z(sum4[2]) );
  CMX2X1 U16 ( .A0(s43[1]), .A1(s44[1]), .S(net107963), .Z(sum4[3]) );
endmodule


module Add_half_3425 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3426 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1713 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3426 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3425 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3427 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3428 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2, n3, n4, n5;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CND2XL U2 ( .A(a), .B(n3), .Z(n4) );
  CND2X1 U3 ( .A(n2), .B(b), .Z(n5) );
  CND2X1 U4 ( .A(n4), .B(n5), .Z(sum) );
  CIVXL U5 ( .A(a), .Z(n2) );
  CIVXL U6 ( .A(b), .Z(n3) );
endmodule


module Add_full_1714 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3428 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3427 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3429 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3430 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2X1 U1 ( .A(n3), .B(n4), .Z(sum) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n1), .B(b), .Z(n4) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1715 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3430 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3429 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_3431 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3432 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net89337, n1, n2, n3, n4;
  assign c_out = net89337;

  CND2X1 U1 ( .A(n1), .B(b), .Z(n4) );
  CND2XL U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVXL U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(net89337) );
endmodule


module Add_full_1716 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3432 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3431 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_429 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1716 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1715 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1714 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1713 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2X1 U3 ( .A(c_out10), .B(n1), .Z(n2) );
  CND2X1 U4 ( .A(n2), .B(n3), .Z(c_out2) );
  CIVX2 U5 ( .A(n4), .Z(n5) );
  CND2X1 U6 ( .A(c_out11), .B(n5), .Z(n3) );
  CIVX1 U7 ( .A(n5), .Z(n1) );
  CMX2X1 U8 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U9 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U10 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n4) );
endmodule


module Add_half_3433 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3434 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1717 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3434 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3433 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3435 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3436 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1718 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3436 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3435 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3437 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3438 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1719 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3438 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3437 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_3439 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3440 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1720 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3440 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3439 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_430 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1720 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1719 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1718 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1717 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n3) );
  CND2X1 U4 ( .A(n5), .B(n6), .Z(c_out2) );
  CND2X1 U5 ( .A(c_out10), .B(n1), .Z(n5) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n3), .Z(n1) );
  CND2IX1 U7 ( .B(n2), .A(n4), .Z(n6) );
  CIVX1 U8 ( .A(c_out11), .Z(n2) );
  CMX2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n4) );
  CMX2XL U10 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U11 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3441 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(n2) );
  CEOXL U3 ( .A(b), .B(n2), .Z(sum) );
  CAN2X1 U4 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3442 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1721 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3442 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3441 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3443 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3444 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1722 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3444 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3443 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3445 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net87260, net106569, net106568, n1;
  assign c_out = net87260;

  CEOX2 U1 ( .A(net106569), .B(b), .Z(sum) );
  CND2X2 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(net87260) );
  CIVXL U4 ( .A(a), .Z(net106568) );
  CIVX1 U5 ( .A(net106568), .Z(net106569) );
endmodule


module Add_half_3446 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88801, n1, n2, n3, n4;
  assign c_out = net88801;

  CIVX2 U1 ( .A(a), .Z(n1) );
  CND2X1 U2 ( .A(a), .B(n2), .Z(n3) );
  CND2X2 U3 ( .A(n1), .B(b), .Z(n4) );
  CND2X2 U4 ( .A(n4), .B(n3), .Z(sum) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(net88801) );
endmodule


module Add_full_1723 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3446 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3445 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVXL U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_3447 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net87261, n1, n2, n3, n4;
  assign c_out = net87261;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CIVX1 U2 ( .A(n2), .Z(net87261) );
  CND2IX1 U3 ( .B(n1), .A(a), .Z(n2) );
  CEOX2 U4 ( .A(n3), .B(b), .Z(sum) );
  CIVX2 U5 ( .A(n4), .Z(n3) );
  CIVXL U6 ( .A(a), .Z(n4) );
endmodule


module Add_half_3448 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88275;
  assign c_out = net88275;

  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(net88275) );
endmodule


module Add_full_1724 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3448 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3447 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_431 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, net76893, n1, n2,
         n3, n4;

  Add_full_1724 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1723 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1722 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1721 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CNIVXL U3 ( .A(net76893), .Z(n1) );
  CIVX2 U4 ( .A(c_out11), .Z(n4) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX1 U6 ( .A(n2), .Z(net76893) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U8 ( .A0(n3), .A1(n4), .S(net76893), .Z(c_out2) );
  CIVX2 U9 ( .A(c_out10), .Z(n3) );
  CMX2XL U10 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
endmodule


module Add_half_3449 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3450 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1725 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3450 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3449 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX2 U1 ( .B(w2), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n1) );
endmodule


module Add_half_3451 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(n2) );
  CEOXL U3 ( .A(b), .B(n2), .Z(sum) );
  CAN2X1 U4 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3452 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1726 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3452 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3451 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3453 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3454 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1727 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3454 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3453 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_3455 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X2 U1 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3456 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1728 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3456 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3455 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_432 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1728 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1727 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1726 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1725 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n2) );
  CMXI2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CIVX2 U5 ( .A(c_out10), .Z(n5) );
  CMX2XL U6 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CMXI2X1 U7 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CMX2XL U8 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U9 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U10 ( .A(c_out11), .Z(n4) );
endmodule


module bit4_108 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, net76936, net76937, net76938,
         net76939, net92795, net92794, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_432 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_431 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_430 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_429 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(c_out401), .A1(c_out400), .S(n1), .Z(n4) );
  CIVX20 U4 ( .A(c_in4), .Z(n1) );
  CIVX1 U5 ( .A(c_out410), .Z(net92795) );
  CMX2X1 U6 ( .A0(c_out401), .A1(c_out400), .S(n3), .Z(n2) );
  CIVX2 U7 ( .A(c_in4), .Z(n3) );
  CMXI2XL U8 ( .A0(n8), .A1(n7), .S(n2), .Z(sum4[3]) );
  CMXI2X1 U9 ( .A0(net92794), .A1(net92795), .S(n4), .Z(c_out4) );
  CMXI2X1 U10 ( .A0(net76938), .A1(net76939), .S(c_in4), .Z(sum4[0]) );
  CMXI2X1 U11 ( .A0(net76936), .A1(net76937), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(c_out411), .Z(net92794) );
  CIVX1 U13 ( .A(s43[0]), .Z(n6) );
  CIVX1 U14 ( .A(s44[1]), .Z(n7) );
  CIVX1 U15 ( .A(s41[1]), .Z(net76936) );
  CIVXL U16 ( .A(s42[1]), .Z(net76937) );
  CIVX2 U17 ( .A(s41[0]), .Z(net76938) );
  CIVX2 U18 ( .A(s42[0]), .Z(net76939) );
  CIVX2 U19 ( .A(s44[0]), .Z(n5) );
  CMXI2X1 U20 ( .A0(n6), .A1(n5), .S(n2), .Z(sum4[2]) );
  CIVX2 U21 ( .A(s43[1]), .Z(n8) );
endmodule


module bit8_27 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, net89764, net89763, net92988,
         net93608, net107934, net76951, net76950, net90088, net93290, net93288,
         net76945, net106472, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_108 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4({b8[3:2], n1, 
        n4}), .c_in4(1'b0) );
  bit4_107 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4({b8[3:2], n1, 
        n4}), .c_in4(1'b1) );
  bit4_106 A83 ( .sum4(s83), .c_out4(c_out810), .a4({a8[7:6], n5, a8[4]}), 
        .b4(b8[7:4]), .c_in4(1'b0) );
  bit4_105 A84 ( .sum4(s84), .c_out4(c_out811), .a4({a8[7:6], n9, a8[4]}), 
        .b4(b8[7:4]), .c_in4(1'b1) );
  CNIVX8 U3 ( .A(b8[0]), .Z(n4) );
  CNIVX4 U4 ( .A(b8[1]), .Z(n1) );
  CMX2X2 U5 ( .A0(s81[3]), .A1(s82[3]), .S(net92988), .Z(sum8[3]) );
  CNIVX3 U6 ( .A(c_in8), .Z(net92988) );
  CIVX2 U7 ( .A(net92988), .Z(net107934) );
  CND2X2 U8 ( .A(net93288), .B(c_out811), .Z(n3) );
  CND2X2 U9 ( .A(n3), .B(net93290), .Z(c_out8) );
  CIVX2 U10 ( .A(net76945), .Z(net93288) );
  CANR2X1 U11 ( .A(n2), .B(c_out800), .C(c_out801), .D(c_in8), .Z(net76945) );
  CND2X1 U12 ( .A(net76945), .B(c_out810), .Z(net93290) );
  CIVX2 U13 ( .A(c_in8), .Z(n2) );
  CMX2X1 U14 ( .A0(s82[2]), .A1(s81[2]), .S(n2), .Z(sum8[2]) );
  CIVXL U15 ( .A(n2), .Z(net106472) );
  CANR2X1 U16 ( .A(c_out800), .B(n2), .C(c_in8), .D(c_out801), .Z(net90088) );
  CANR2XL U17 ( .A(net107934), .B(c_out800), .C(net106472), .D(c_out801), .Z(
        net89763) );
  CANR2X1 U18 ( .A(c_out800), .B(net93608), .C(c_in8), .D(c_out801), .Z(
        net89764) );
  CMXI2X1 U19 ( .A0(net76950), .A1(net76951), .S(net90088), .Z(sum8[4]) );
  CIVX2 U20 ( .A(s83[0]), .Z(net76951) );
  CIVX2 U21 ( .A(s84[0]), .Z(net76950) );
  CIVX1 U22 ( .A(s83[2]), .Z(n14) );
  CIVX3 U23 ( .A(n8), .Z(n5) );
  CIVX3 U24 ( .A(n8), .Z(n9) );
  CND2X2 U25 ( .A(s81[1]), .B(net107934), .Z(n6) );
  CND2X1 U26 ( .A(s82[1]), .B(net92988), .Z(n7) );
  CND2X4 U27 ( .A(n6), .B(n7), .Z(sum8[1]) );
  CIVXL U28 ( .A(c_in8), .Z(net93608) );
  CIVX1 U29 ( .A(s84[2]), .Z(n15) );
  CMX2X2 U30 ( .A0(s84[3]), .A1(s83[3]), .S(net89763), .Z(sum8[7]) );
  CIVX2 U31 ( .A(a8[5]), .Z(n8) );
  CMXI2X1 U32 ( .A0(n11), .A1(n10), .S(c_in8), .Z(sum8[0]) );
  CMXI2X1 U33 ( .A0(n13), .A1(n12), .S(net89764), .Z(sum8[5]) );
  CMXI2X1 U34 ( .A0(n15), .A1(n14), .S(net89764), .Z(sum8[6]) );
  CIVX2 U35 ( .A(s81[0]), .Z(n11) );
  CIVX2 U36 ( .A(s82[0]), .Z(n10) );
  CIVX2 U37 ( .A(s84[1]), .Z(n13) );
  CIVX2 U38 ( .A(s83[1]), .Z(n12) );
endmodule


module Add_half_3457 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3458 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1729 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3458 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3457 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3459 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3460 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1730 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3460 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3459 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3461 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3462 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1731 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3462 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3461 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3463 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3464 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1732 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3464 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3463 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_433 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_1732 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1731 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1730 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1729 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CIVX2 U4 ( .A(c_in2), .Z(n2) );
  CMX2X1 U5 ( .A0(c_out11), .A1(c_out10), .S(n3), .Z(c_out2) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n3) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3465 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3466 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1733 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3466 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3465 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3467 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3468 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1734 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3468 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3467 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3469 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3470 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1735 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3470 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3469 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3471 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3472 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1736 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3472 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3471 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_434 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1736 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1735 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1734 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1733 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2X1 U4 ( .A0(c_out11), .A1(c_out10), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CIVX2 U7 ( .A(s1), .Z(n4) );
  CIVX2 U8 ( .A(s2), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3473 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3474 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1737 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3474 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3473 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3475 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3476 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1738 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3476 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3475 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3477 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CAN2X2 U1 ( .A(b), .B(a), .Z(c_out) );
  CIVXL U2 ( .A(a), .Z(n1) );
  CIVX1 U3 ( .A(n1), .Z(n2) );
  CEOXL U4 ( .A(n2), .B(b), .Z(sum) );
endmodule


module Add_half_3478 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1739 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3478 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3477 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3479 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3480 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1740 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3480 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3479 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_435 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, net77054,
         net77055, net91751, n1, n2, n3, n4, n5, n6;

  Add_full_1740 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1739 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1738 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1737 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CANR2X2 U4 ( .A(n4), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n1) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CANR2XL U6 ( .A(n4), .B(c_out00), .C(c_in2), .D(c_out01), .Z(net91751) );
  CIVX2 U7 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(net77054), .A1(net77055), .S(c_in2), .Z(sum2[0]) );
  CIVX1 U10 ( .A(s2), .Z(net77055) );
  CIVX1 U11 ( .A(s1), .Z(net77054) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
  CIVX2 U13 ( .A(s3), .Z(n5) );
  CMXI2X1 U14 ( .A0(n6), .A1(n5), .S(net91751), .Z(sum2[1]) );
endmodule


module Add_half_3481 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3482 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1741 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3482 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3481 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3483 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3484 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1742 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3484 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3483 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3485 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3486 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   net88512;
  assign c_out = net88512;

  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(net88512) );
endmodule


module Add_full_1743 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3486 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3485 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3487 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n3;

  CNIVX1 U1 ( .A(a), .Z(n1) );
  CENX1 U2 ( .A(n3), .B(n1), .Z(sum) );
  CAN2X1 U3 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U4 ( .A(b), .Z(n3) );
endmodule


module Add_half_3488 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1744 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3488 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3487 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_436 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, net92672,
         net77089, net77088, n1, n2, n3, n4;

  Add_full_1744 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1743 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1742 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1741 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CND2X2 U4 ( .A(n1), .B(c_out00), .Z(n3) );
  CND2IX2 U5 ( .B(n1), .A(c_out01), .Z(n4) );
  CND2X2 U6 ( .A(n3), .B(n4), .Z(n2) );
  CMXI2X1 U7 ( .A0(net77089), .A1(net77088), .S(n2), .Z(c_out2) );
  CMXI2XL U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(net92672) );
  CMX2XL U9 ( .A0(s4), .A1(s3), .S(net92672), .Z(sum2[1]) );
  CMX2X1 U10 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(c_out10), .Z(net77089) );
  CIVX2 U12 ( .A(c_out11), .Z(net77088) );
endmodule


module bit4_109 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, net91766, net77101, net77100,
         n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_436 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_435 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_434 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_433 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n3) );
  CNIVX1 U4 ( .A(net91766), .Z(n1) );
  CMXI2X1 U5 ( .A0(net77100), .A1(net77101), .S(n3), .Z(c_out4) );
  CIVX2 U6 ( .A(c_in4), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out401), .A1(c_out400), .S(n2), .Z(net91766) );
  CMXI2X1 U8 ( .A0(n5), .A1(n4), .S(n1), .Z(sum4[3]) );
  CIVX1 U9 ( .A(c_out410), .Z(net77101) );
  CIVX1 U10 ( .A(c_out411), .Z(net77100) );
  CMX2X1 U11 ( .A0(s44[0]), .A1(s43[0]), .S(net91766), .Z(sum4[2]) );
  CMX2X1 U12 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U13 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX1 U14 ( .A(s44[1]), .Z(n5) );
  CIVX2 U15 ( .A(s43[1]), .Z(n4) );
endmodule


module Add_half_3489 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3490 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1745 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3490 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3489 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3491 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3492 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1746 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3492 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3491 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3493 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3494 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1747 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3494 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3493 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3495 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3496 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1748 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3496 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3495 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_437 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1748 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1747 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1746 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1745 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2X1 U4 ( .A0(c_out11), .A1(c_out10), .S(n2), .Z(c_out2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module Add_half_3497 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3498 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1749 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3498 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3497 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3499 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3500 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1750 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3500 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3499 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3501 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3502 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1751 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3502 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3501 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3503 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3504 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1752 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3504 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3503 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CNR2X1 U2 ( .A(w3), .B(w2), .Z(n1) );
endmodule


module bit2_438 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_1752 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1751 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1750 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1749 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2XL U4 ( .A0(n3), .A1(n2), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(s3), .Z(n3) );
  CIVX2 U8 ( .A(s4), .Z(n2) );
endmodule


module Add_half_3505 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3506 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1753 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3506 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3505 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3507 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3508 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1754 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3508 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3507 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3509 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3510 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1755 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3510 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3509 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3511 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n4;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(n2) );
  CENXL U3 ( .A(n4), .B(n2), .Z(sum) );
  CAN2X1 U4 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U5 ( .A(b), .Z(n4) );
endmodule


module Add_half_3512 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4, n5;

  CND2XL U1 ( .A(n2), .B(a), .Z(n5) );
  CIVXL U2 ( .A(n3), .Z(n1) );
  CIVX1 U3 ( .A(a), .Z(n3) );
  CND2X1 U4 ( .A(b), .B(n3), .Z(n4) );
  CND2X1 U5 ( .A(n4), .B(n5), .Z(sum) );
  CIVX1 U6 ( .A(b), .Z(n2) );
  CAN2XL U7 ( .A(b), .B(n1), .Z(c_out) );
endmodule


module Add_full_1756 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3512 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3511 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_439 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1756 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1755 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1754 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1753 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2XL U3 ( .A(n2), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n1) );
  CANR2X2 U4 ( .A(c_out00), .B(n2), .C(c_in2), .D(c_out01), .Z(n5) );
  CMX2XL U5 ( .A0(s4), .A1(s3), .S(n1), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out11), .Z(n4) );
  CIVX2 U8 ( .A(c_out10), .Z(n3) );
  CIVX2 U9 ( .A(c_in2), .Z(n2) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(n5), .Z(c_out2) );
endmodule


module Add_half_3513 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3514 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1757 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3514 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3513 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3515 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3516 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1758 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3516 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3515 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3517 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOX1 U1 ( .A(b), .B(n1), .Z(sum) );
  CNIVXL U2 ( .A(a), .Z(n1) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3518 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3;

  CND2IXL U1 ( .B(b), .A(a), .Z(n3) );
  CND2X2 U2 ( .A(b), .B(n1), .Z(n2) );
  CND2X2 U3 ( .A(n2), .B(n3), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CAN2XL U5 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1759 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3518 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3517 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3519 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3520 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1760 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3520 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3519 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_440 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1760 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1759 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1758 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1757 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X2 U3 ( .A(n1), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n4) );
  CMX2XL U4 ( .A0(s4), .A1(s3), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out11), .Z(n3) );
  CIVX2 U7 ( .A(c_out10), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_110 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_440 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_439 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_438 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_437 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(n10), .Z(n1) );
  CMX2X1 U4 ( .A0(s42[0]), .A1(s41[0]), .S(n5), .Z(sum4[0]) );
  CMXI2X1 U5 ( .A0(n9), .A1(n8), .S(n4), .Z(sum4[2]) );
  CMX2XL U6 ( .A0(s44[1]), .A1(s43[1]), .S(n4), .Z(sum4[3]) );
  CND2X2 U7 ( .A(n2), .B(n3), .Z(c_out4) );
  CND2X2 U8 ( .A(c_out411), .B(n1), .Z(n2) );
  CND2X1 U9 ( .A(c_out410), .B(n10), .Z(n3) );
  CANR2X1 U10 ( .A(c_out400), .B(n5), .C(c_in4), .D(c_out401), .Z(n4) );
  CANR2X1 U11 ( .A(c_out400), .B(n5), .C(c_out401), .D(c_in4), .Z(n10) );
  CIVX2 U12 ( .A(c_in4), .Z(n5) );
  CIVX2 U13 ( .A(s41[1]), .Z(n7) );
  CIVX2 U14 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U15 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U16 ( .A(s44[0]), .Z(n9) );
  CIVX2 U17 ( .A(s43[0]), .Z(n8) );
endmodule


module Add_half_3521 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3522 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1761 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3522 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3521 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3523 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3524 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1762 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3524 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3523 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3525 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n4;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(n2) );
  CENXL U3 ( .A(n4), .B(n2), .Z(sum) );
  CAN2X1 U4 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U5 ( .A(b), .Z(n4) );
endmodule


module Add_half_3526 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1763 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3526 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3525 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3527 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_3528 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1764 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3528 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3527 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_441 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1764 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1763 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1762 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1761 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s3), .Z(n4) );
  CIVX2 U9 ( .A(s4), .Z(n3) );
endmodule


module Add_half_3529 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_3530 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX2 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1765 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3530 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3529 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3531 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
  CIVX2 U4 ( .A(b), .Z(n2) );
endmodule


module Add_half_3532 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_full_1766 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3532 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3531 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3533 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3534 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1767 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3534 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3533 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3535 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X2 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3536 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1768 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3536 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3535 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_442 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1768 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1767 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1766 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1765 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_3537 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3538 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1769 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3538 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3537 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3539 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3540 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1770 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3540 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3539 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3541 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3542 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1771 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3542 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3541 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3543 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CEOXL U2 ( .A(n1), .B(b), .Z(sum) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3544 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1772 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3544 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3543 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_443 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1772 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1771 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1770 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1769 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CIVX1 U5 ( .A(n2), .Z(n5) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n4) );
  CIVX2 U8 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n5), .Z(c_out2) );
  CIVX2 U10 ( .A(s3), .Z(n7) );
  CIVX2 U11 ( .A(s4), .Z(n6) );
  CMXI2X1 U12 ( .A0(n7), .A1(n6), .S(n5), .Z(sum2[1]) );
endmodule


module Add_half_3545 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3546 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX1 U1 ( .A(a), .B(n1), .Z(sum) );
  CIVX2 U2 ( .A(b), .Z(n1) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1773 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3546 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3545 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3547 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3548 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1774 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3548 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3547 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3549 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3550 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1775 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3550 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3549 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3551 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3552 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1776 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3552 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3551 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_444 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1776 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1775 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1774 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1773 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(c_out10), .Z(n3) );
  CIVX1 U4 ( .A(n1), .Z(n6) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX1 U6 ( .A(s1), .Z(n5) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module bit4_111 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_444 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_443 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_442 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_441 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2X1 U4 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2XL U5 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U7 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX1 U8 ( .A(c_out410), .Z(n3) );
  CIVX2 U9 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module Add_half_3553 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3554 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_full_1777 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3554 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3553 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3555 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_3556 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX2 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1778 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3556 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3555 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3557 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3558 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2, n3, n4;

  CND2XL U1 ( .A(a), .B(n2), .Z(n3) );
  CND2X2 U2 ( .A(n1), .B(b), .Z(n4) );
  CND2X2 U3 ( .A(n3), .B(n4), .Z(sum) );
  CIVX1 U4 ( .A(a), .Z(n1) );
  CIVXL U5 ( .A(b), .Z(n2) );
  CAN2XL U6 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1779 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3558 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3557 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3559 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X2 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3560 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1780 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3560 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3559 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_445 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1780 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1779 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1778 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1777 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(c_out11), .Z(n4) );
  CMX2X1 U4 ( .A0(s3), .A1(s4), .S(n8), .Z(sum2[1]) );
  CIVX1 U5 ( .A(s2), .Z(n6) );
  CIVX1 U6 ( .A(s1), .Z(n7) );
  CIVXL U7 ( .A(n2), .Z(n1) );
  CIVX2 U8 ( .A(n3), .Z(n2) );
  CIVXL U9 ( .A(n1), .Z(n8) );
  CIVX2 U10 ( .A(c_out10), .Z(n5) );
  CMXI2X1 U11 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n3) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(n2), .Z(c_out2) );
  CMXI2X1 U13 ( .A0(n7), .A1(n6), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_3561 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_3562 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CIVX2 U1 ( .A(b), .Z(n2) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_full_1781 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3562 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3561 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_3563 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_3564 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_full_1782 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3564 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3563 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_3565 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3566 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1783 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3566 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3565 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3567 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3568 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1784 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3568 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3567 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_446 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1784 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1783 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1782 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1781 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2X1 U3 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CIVX2 U4 ( .A(c_in2), .Z(n2) );
  CMX2XL U5 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n3) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(c_out10), .Z(n5) );
  CIVX2 U10 ( .A(c_out11), .Z(n4) );
endmodule


module Add_half_3569 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3570 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVXL U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1785 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3570 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3569 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3571 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3572 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1786 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3572 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3571 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3573 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3574 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1787 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3574 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3573 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3575 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3576 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1788 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3576 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3575 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_447 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1788 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1787 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1786 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1785 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX1 U4 ( .A(c_out10), .Z(n3) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_3577 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3578 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVXL U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1789 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3578 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3577 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3579 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3580 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVXL U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1790 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3580 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3579 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3581 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3582 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1791 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3582 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3581 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3583 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3584 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1792 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3584 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3583 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_448 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1792 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1791 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1790 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1789 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(c_out10), .Z(n3) );
  CIVX1 U4 ( .A(c_out11), .Z(n2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_112 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_448 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_447 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_446 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_445 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(n4), .A1(n3), .S(n1), .Z(c_out4) );
  CMX2X1 U4 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U5 ( .A(s44[1]), .Z(n12) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CIVX1 U7 ( .A(c_out411), .Z(n3) );
  CIVX1 U8 ( .A(c_out410), .Z(n4) );
  CIVX1 U9 ( .A(s41[1]), .Z(n8) );
  CIVX1 U10 ( .A(s41[0]), .Z(n6) );
  CIVX2 U11 ( .A(n2), .Z(n11) );
  CIVX2 U12 ( .A(s42[0]), .Z(n5) );
  CMXI2X1 U13 ( .A0(n6), .A1(n5), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U14 ( .A(s42[1]), .Z(n7) );
  CMXI2X1 U15 ( .A0(n8), .A1(n7), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U16 ( .A(s43[0]), .Z(n10) );
  CIVX2 U17 ( .A(s44[0]), .Z(n9) );
  CMXI2X1 U18 ( .A0(n10), .A1(n9), .S(n11), .Z(sum4[2]) );
  CIVX2 U19 ( .A(s43[1]), .Z(n13) );
  CMXI2X1 U20 ( .A0(n13), .A1(n12), .S(n11), .Z(sum4[3]) );
endmodule


module bit8_28 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   n26, c_out800, c_out801, c_out810, c_out811, net77525, net77542,
         net77540, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_112 A81 ( .sum4(s81), .c_out4(c_out800), .a4({n11, a8[2:0]}), .b4({
        b8[3], n12, b8[1:0]}), .c_in4(1'b0) );
  bit4_111 A82 ( .sum4(s82), .c_out4(c_out801), .a4({n11, a8[2:0]}), .b4({
        b8[3], n12, b8[1:0]}), .c_in4(1'b1) );
  bit4_110 A83 ( .sum4(s83), .c_out4(c_out810), .a4({a8[7:5], n17}), .b4({
        b8[7:5], n9}), .c_in4(1'b0) );
  bit4_109 A84 ( .sum4(s84), .c_out4(c_out811), .a4({a8[7:5], n3}), .b4({
        b8[7:5], n2}), .c_in4(1'b1) );
  CIVDX2 U3 ( .A(b8[4]), .Z0(n1), .Z1(n2) );
  CMX2X2 U4 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CNIVX4 U5 ( .A(b8[2]), .Z(n12) );
  CMXI2X2 U6 ( .A0(n19), .A1(n18), .S(c_in8), .Z(sum8[0]) );
  CMXI2X2 U7 ( .A0(n21), .A1(n20), .S(c_in8), .Z(sum8[1]) );
  CIVX4 U8 ( .A(n1), .Z(n9) );
  CIVX4 U9 ( .A(n16), .Z(n3) );
  CIVX3 U10 ( .A(n16), .Z(n17) );
  CIVXL U11 ( .A(net77525), .Z(n4) );
  CIVX1 U12 ( .A(n4), .Z(n5) );
  CMX2X1 U13 ( .A0(s83[3]), .A1(s84[3]), .S(n5), .Z(n26) );
  CND2XL U14 ( .A(s83[2]), .B(n6), .Z(n7) );
  CND2XL U15 ( .A(s84[2]), .B(net77525), .Z(n8) );
  CND2X1 U16 ( .A(n7), .B(n8), .Z(sum8[6]) );
  CIVXL U17 ( .A(net77525), .Z(n6) );
  CIVX4 U18 ( .A(a8[3]), .Z(n10) );
  CIVX8 U19 ( .A(n10), .Z(n11) );
  CIVX1 U20 ( .A(s83[0]), .Z(n25) );
  CND2X4 U21 ( .A(net77540), .B(n13), .Z(c_out8) );
  CND2IX2 U22 ( .B(n14), .A(c_out811), .Z(n13) );
  CMXI2XL U23 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n14) );
  CND2IX2 U24 ( .B(net77525), .A(c_out810), .Z(net77540) );
  CIVX2 U25 ( .A(net77542), .Z(net77525) );
  CMXI2X1 U26 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(net77542) );
  CNIVX4 U27 ( .A(n26), .Z(sum8[7]) );
  CMX2X2 U28 ( .A0(s83[1]), .A1(s84[1]), .S(net77525), .Z(sum8[5]) );
  CIVX2 U29 ( .A(a8[4]), .Z(n16) );
  CMXI2X1 U30 ( .A0(n25), .A1(n24), .S(net77525), .Z(sum8[4]) );
  CIVX1 U31 ( .A(s81[1]), .Z(n21) );
  CIVX1 U32 ( .A(s82[1]), .Z(n20) );
  CIVX1 U33 ( .A(s82[0]), .Z(n18) );
  CIVX1 U34 ( .A(s81[0]), .Z(n19) );
  CIVX1 U35 ( .A(s82[2]), .Z(n22) );
  CIVX1 U36 ( .A(s81[2]), .Z(n23) );
  CMXI2X1 U37 ( .A0(n23), .A1(n22), .S(c_in8), .Z(sum8[2]) );
  CIVX2 U38 ( .A(s84[0]), .Z(n24) );
endmodule


module bit32_7 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   n3, c1, c2, c3, n1;

  bit8_28 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8({a32[7:2], n1, a32[0]}), 
        .b8(b32[7:0]), .c_in8(c_in32) );
  bit8_27 A322 ( .sum8({sum32[15:11], n3, sum32[9:8]}), .c_out8(c2), .a8(
        a32[15:8]), .b8(b32[15:8]), .c_in8(c1) );
  bit8_26 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8(a32[23:16]), .b8(
        b32[23:16]), .c_in8(c2) );
  bit8_25 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8(a32[31:24]), .b8(
        b32[31:24]), .c_in8(c3) );
  CNIVX4 U1 ( .A(a32[1]), .Z(n1) );
  CNIVX4 U2 ( .A(n3), .Z(sum32[10]) );
endmodule


module Add_half_3585 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3586 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1793 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3586 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3585 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3587 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3588 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1794 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3588 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3587 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3589 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3590 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1795 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3590 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3589 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3591 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3592 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1796 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3592 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3591 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_449 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1796 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1795 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1794 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1793 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3593 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3594 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1797 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3594 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3593 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3595 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3596 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1798 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3596 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3595 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3597 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3598 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1799 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3598 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3597 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3599 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3600 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1800 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3600 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3599 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_450 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1800 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1799 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1798 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1797 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3601 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3602 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1801 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3602 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3601 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3603 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3604 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1802 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3604 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3603 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3605 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3606 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1803 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3606 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3605 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3607 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3608 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1804 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3608 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3607 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_451 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1804 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1803 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1802 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1801 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3609 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3610 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1805 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3610 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3609 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3611 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3612 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1806 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3612 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3611 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3613 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3614 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1807 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3614 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3613 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3615 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3616 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1808 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3616 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3615 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_452 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1808 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1807 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1806 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1805 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_113 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_452 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_451 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_450 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_449 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_3617 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3618 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1809 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3618 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3617 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3619 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3620 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1810 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3620 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3619 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3621 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3622 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1811 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3622 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3621 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3623 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3624 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1812 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3624 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3623 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_453 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1812 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1811 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1810 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1809 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3625 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3626 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1813 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3626 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3625 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3627 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3628 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1814 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3628 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3627 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3629 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3630 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1815 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3630 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3629 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3631 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3632 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1816 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3632 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3631 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_454 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1816 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1815 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1814 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1813 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3633 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3634 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1817 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3634 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3633 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3635 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3636 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1818 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3636 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3635 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3637 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3638 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1819 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3638 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3637 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3639 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3640 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1820 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3640 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3639 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_455 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1820 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1819 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1818 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1817 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3641 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3642 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1821 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3642 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3641 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3643 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3644 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1822 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3644 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3643 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3645 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3646 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1823 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3646 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3645 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3647 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3648 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1824 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3648 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3647 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_456 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1824 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1823 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1822 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1821 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_114 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_456 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_455 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_454 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_453 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_3649 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3650 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1825 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3650 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3649 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3651 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3652 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1826 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3652 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3651 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3653 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3654 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1827 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3654 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3653 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3655 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3656 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1828 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3656 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3655 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_457 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1828 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1827 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1826 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1825 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3657 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3658 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1829 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3658 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3657 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3659 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3660 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1830 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3660 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3659 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3661 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3662 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1831 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3662 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3661 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3663 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3664 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1832 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3664 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3663 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_458 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1832 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1831 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1830 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1829 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3665 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3666 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1833 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3666 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3665 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3667 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3668 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1834 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3668 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3667 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3669 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3670 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1835 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3670 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3669 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3671 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3672 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1836 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3672 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3671 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_459 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1836 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1835 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1834 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1833 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CAOR2XL U3 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CANR2X1 U7 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3673 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3674 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1837 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3674 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3673 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3675 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3676 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1838 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3676 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3675 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3677 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3678 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1839 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3678 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3677 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3679 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3680 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1840 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3680 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3679 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_460 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1840 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1839 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1838 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1837 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_115 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_460 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_459 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_458 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_457 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
endmodule


module Add_half_3681 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3682 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1841 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3682 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3681 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3683 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3684 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1842 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3684 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3683 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3685 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3686 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1843 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3686 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3685 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3687 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3688 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1844 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3688 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3687 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_461 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1844 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1843 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1842 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1841 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CAOR2XL U3 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CANR2X1 U6 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3689 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3690 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1845 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3690 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3689 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3691 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3692 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1846 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3692 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3691 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3693 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3694 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1847 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3694 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3693 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3695 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3696 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1848 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3696 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3695 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_462 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1848 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1847 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1846 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1845 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3697 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3698 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1849 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3698 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3697 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3699 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3700 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1850 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3700 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3699 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3701 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3702 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1851 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3702 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3701 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3703 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3704 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1852 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3704 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3703 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_463 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1852 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1851 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1850 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1849 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CAOR2XL U3 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CANR2X1 U6 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3705 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3706 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1853 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3706 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3705 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3707 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3708 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1854 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3708 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3707 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3709 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3710 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1855 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3710 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3709 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3711 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3712 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1856 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3712 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3711 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_464 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1856 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1855 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1854 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1853 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_116 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_464 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_463 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_462 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_461 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2XL U3 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U10 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_29 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_116 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_115 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_114 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_113 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out8) );
  CMX2X1 U4 ( .A0(s83[3]), .A1(s84[3]), .S(n1), .Z(sum8[7]) );
  CMX2X1 U5 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CMX2X1 U6 ( .A0(s83[2]), .A1(s84[2]), .S(n1), .Z(sum8[6]) );
  CMX2X1 U7 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CIVX1 U8 ( .A(s82[0]), .Z(n4) );
  CMX2X1 U9 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2X1 U10 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2X1 U11 ( .A0(s83[0]), .A1(s84[0]), .S(n1), .Z(sum8[4]) );
  CMX2X1 U12 ( .A0(s83[1]), .A1(s84[1]), .S(n1), .Z(sum8[5]) );
  CIVX2 U13 ( .A(c_out810), .Z(n3) );
  CIVX2 U14 ( .A(c_out811), .Z(n2) );
  CIVX2 U15 ( .A(s81[0]), .Z(n5) );
  CMXI2X1 U16 ( .A0(n5), .A1(n4), .S(c_in8), .Z(sum8[0]) );
endmodule


module Add_half_3713 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3714 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1857 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3714 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3713 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3715 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3716 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1858 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3716 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3715 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3717 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3718 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1859 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3718 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3717 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3719 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3720 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1860 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3720 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3719 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_465 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1860 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1859 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1858 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1857 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_3721 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3722 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1861 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3722 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3721 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3723 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3724 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1862 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3724 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3723 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3725 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3726 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1863 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3726 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3725 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3727 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3728 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1864 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3728 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3727 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_466 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1864 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1863 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1862 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1861 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CIVXL U3 ( .A(s3), .Z(n4) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_3729 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3730 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1865 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3730 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3729 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3731 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3732 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1866 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3732 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3731 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3733 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3734 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1867 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3734 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3733 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3735 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3736 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1868 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3736 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3735 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_467 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1868 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1867 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1866 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1865 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_3737 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_3738 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1869 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3738 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3737 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3739 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3740 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1870 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3740 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3739 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3741 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3742 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1871 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3742 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3741 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3743 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3744 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1872 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3744 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3743 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_468 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_1872 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1871 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1870 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1869 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVXL U3 ( .A(s3), .Z(n6) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module bit4_117 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_468 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_467 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_466 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_465 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n3), .Z(sum4[0]) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n2), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n2), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(c_out410), .A1(c_out411), .S(n2), .Z(c_out4) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMXI2X1 U7 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n2) );
  CIVX2 U10 ( .A(c_in4), .Z(n3) );
endmodule


module Add_half_3745 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3746 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1873 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3746 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3745 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3747 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3748 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1874 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3748 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3747 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3749 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3750 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1875 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3750 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3749 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3751 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3752 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1876 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3752 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3751 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_469 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1876 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1875 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1874 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1873 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_3753 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3754 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1877 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3754 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3753 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3755 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3756 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1878 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3756 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3755 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3757 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3758 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1879 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3758 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3757 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3759 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3760 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1880 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3760 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3759 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_470 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1880 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1879 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1878 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1877 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_3761 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3762 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1881 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3762 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3761 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3763 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3764 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1882 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3764 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3763 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3765 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3766 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1883 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3766 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3765 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3767 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3768 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1884 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3768 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3767 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_471 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1884 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1883 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1882 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1881 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_3769 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3770 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1885 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3770 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3769 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3771 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3772 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1886 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3772 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3771 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3773 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3774 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1887 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3774 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3773 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3775 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3776 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1888 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3776 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3775 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_472 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1888 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1887 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1886 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1885 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module bit4_118 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_472 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_471 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_470 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_469 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n11), .Z(sum4[0]) );
  CIVX2 U3 ( .A(c_out410), .Z(n3) );
  CIVX2 U4 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n8) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U8 ( .A(s41[1]), .Z(n5) );
  CIVX2 U10 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(s43[0]), .Z(n7) );
  CIVX2 U13 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX2 U15 ( .A(s43[1]), .Z(n10) );
  CIVX2 U16 ( .A(s44[1]), .Z(n9) );
  CMXI2X1 U17 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
  CIVX2 U18 ( .A(c_in4), .Z(n11) );
endmodule


module Add_half_3777 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3778 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1889 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3778 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3777 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3779 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3780 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1890 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3780 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3779 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3781 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3782 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1891 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3782 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3781 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3783 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3784 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1892 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3784 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3783 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_473 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_1892 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1891 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1890 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1889 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_3785 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3786 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1893 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3786 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3785 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3787 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3788 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1894 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3788 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3787 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3789 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3790 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1895 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3790 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3789 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3791 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3792 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1896 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3792 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3791 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_474 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_1896 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1895 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1894 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1893 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_3793 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3794 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1897 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3794 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3793 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3795 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3796 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1898 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3796 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3795 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3797 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3798 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1899 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3798 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3797 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3799 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3800 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1900 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3800 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3799 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_475 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1900 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1899 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1898 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1897 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_3801 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3802 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1901 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3802 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3801 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3803 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3804 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1902 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3804 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3803 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3805 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3806 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1903 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3806 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3805 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3807 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3808 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1904 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3808 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3807 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_476 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_1904 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1903 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1902 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1901 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_119 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_476 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_475 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_474 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_473 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(c_out410), .Z(n3) );
  CIVX2 U4 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n10) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n10), .Z(c_out4) );
  CIVX2 U8 ( .A(s41[0]), .Z(n5) );
  CIVX2 U9 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U11 ( .A(s41[1]), .Z(n7) );
  CIVX2 U12 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U13 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n9) );
  CIVX2 U15 ( .A(s44[0]), .Z(n8) );
  CMXI2X1 U16 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CIVX2 U17 ( .A(s43[1]), .Z(n12) );
  CIVX2 U18 ( .A(s44[1]), .Z(n11) );
  CMXI2X1 U19 ( .A0(n12), .A1(n11), .S(n10), .Z(sum4[3]) );
endmodule


module Add_half_3809 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3810 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1905 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3810 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3809 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3811 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3812 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1906 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3812 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3811 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3813 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3814 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1907 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3814 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3813 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3815 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3816 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1908 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3816 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3815 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_477 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1908 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1907 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1906 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1905 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CIVXL U3 ( .A(s3), .Z(n4) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_3817 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3818 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1909 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3818 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3817 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3819 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3820 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1910 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3820 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3819 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3821 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3822 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1911 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3822 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3821 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3823 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3824 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1912 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3824 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3823 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_478 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_1912 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1911 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1910 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1909 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(n1), .Z(n2) );
  CIVX2 U6 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_3825 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3826 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1913 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3826 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3825 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3827 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3828 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1914 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3828 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3827 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3829 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3830 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1915 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3830 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3829 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3831 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3832 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1916 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3832 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3831 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_479 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1916 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1915 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1914 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1913 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(s3), .Z(n8) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_3833 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3834 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1917 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3834 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3833 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3835 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3836 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1918 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3836 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3835 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3837 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3838 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1919 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3838 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3837 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3839 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_3840 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1920 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3840 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3839 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_480 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1920 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1919 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1918 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1917 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module bit4_120 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_480 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_479 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_478 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_477 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module bit8_30 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_120 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_119 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_118 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_117 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X1 U3 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2XL U4 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2X1 U5 ( .A0(s83[2]), .A1(s84[2]), .S(n2), .Z(sum8[6]) );
  CMX2X1 U6 ( .A0(s81[0]), .A1(s82[0]), .S(c_in8), .Z(sum8[0]) );
  CMX2X2 U7 ( .A0(s83[0]), .A1(s84[0]), .S(n2), .Z(sum8[4]) );
  CMX2X1 U8 ( .A0(c_out810), .A1(c_out811), .S(n2), .Z(c_out8) );
  CIVX2 U9 ( .A(n1), .Z(n2) );
  CMX2X1 U10 ( .A0(s83[3]), .A1(s84[3]), .S(n2), .Z(sum8[7]) );
  CMX2X1 U11 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2X1 U12 ( .A0(s83[1]), .A1(s84[1]), .S(n2), .Z(sum8[5]) );
  CMXI2X1 U13 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
endmodule


module Add_half_3841 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3842 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1921 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3842 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3841 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3843 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3844 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1922 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3844 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3843 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3845 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3846 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1923 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3846 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3845 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_3847 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3848 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1924 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3848 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3847 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_481 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_1924 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1923 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1922 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1921 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(s4), .Z(n7) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s3), .Z(n8) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_3849 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3850 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1925 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3850 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3849 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3851 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3852 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1926 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3852 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3851 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3853 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_3854 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1927 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3854 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3853 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3855 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3856 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1928 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_3856 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3855 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_482 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_1928 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1927 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1926 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1925 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_3857 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3858 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1929 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3858 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3857 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3859 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3860 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1930 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3860 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3859 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3861 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3862 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1931 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3862 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3861 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3863 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3864 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1932 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3864 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3863 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_483 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1932 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1931 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1930 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1929 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3865 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3866 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1933 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3866 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3865 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3867 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3868 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1934 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3868 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3867 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3869 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3870 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1935 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3870 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3869 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3871 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3872 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1936 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3872 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3871 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_484 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1936 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1935 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1934 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1933 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_121 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_484 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_483 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_482 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_481 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMX2X1 U4 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CMX2X1 U5 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U6 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_3873 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3874 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1937 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3874 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3873 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3875 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3876 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1938 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3876 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3875 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3877 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3878 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1939 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3878 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3877 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_3879 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3880 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1940 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3880 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3879 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_485 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1940 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1939 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1938 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1937 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_3881 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3882 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1941 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3882 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3881 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3883 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3884 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_1942 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3884 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3883 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_3885 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3886 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1943 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3886 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3885 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_3887 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_3888 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_1944 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_3888 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3887 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_486 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_1944 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1943 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1942 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1941 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_3889 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3890 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1945 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3890 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3889 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3891 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3892 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1946 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3892 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3891 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3893 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3894 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1947 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3894 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3893 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3895 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3896 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1948 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3896 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3895 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_487 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1948 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1947 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1946 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1945 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3897 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3898 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1949 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3898 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3897 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3899 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3900 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1950 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3900 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3899 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3901 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3902 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1951 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3902 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3901 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3903 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3904 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1952 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3904 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3903 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_488 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1952 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1951 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1950 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1949 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_122 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_488 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_487 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_486 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_485 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n8), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n8), .Z(sum4[0]) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U4 ( .A(c_out410), .Z(n3) );
  CIVX2 U5 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U6 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out4) );
  CIVX2 U7 ( .A(s43[0]), .Z(n5) );
  CIVX2 U10 ( .A(s44[0]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(n1), .Z(sum4[2]) );
  CIVX2 U12 ( .A(s43[1]), .Z(n7) );
  CIVX2 U13 ( .A(s44[1]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n1), .Z(sum4[3]) );
  CIVX2 U15 ( .A(c_in4), .Z(n8) );
endmodule


module Add_half_3905 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3906 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1953 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3906 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3905 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3907 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3908 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1954 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3908 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3907 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3909 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3910 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1955 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3910 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3909 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3911 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3912 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1956 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3912 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3911 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_489 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1956 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1955 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1954 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1953 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3913 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3914 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1957 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3914 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3913 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3915 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3916 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1958 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3916 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3915 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3917 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3918 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1959 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3918 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3917 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3919 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3920 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1960 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3920 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3919 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_490 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1960 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1959 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1958 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1957 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3921 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3922 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1961 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3922 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3921 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3923 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3924 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1962 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3924 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3923 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3925 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3926 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1963 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3926 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3925 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3927 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3928 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1964 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3928 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3927 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_491 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1964 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1963 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1962 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1961 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3929 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3930 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1965 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3930 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3929 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3931 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3932 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1966 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3932 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3931 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3933 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3934 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1967 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3934 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3933 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3935 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3936 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1968 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3936 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3935 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_492 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1968 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1967 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1966 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1965 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_123 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_492 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_491 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_490 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_489 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_3937 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3938 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1969 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3938 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3937 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3939 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3940 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1970 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3940 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3939 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3941 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3942 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1971 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3942 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3941 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3943 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3944 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1972 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3944 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3943 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_493 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1972 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1971 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1970 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1969 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3945 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3946 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1973 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3946 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3945 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3947 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3948 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1974 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3948 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3947 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3949 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3950 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1975 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3950 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3949 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3951 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3952 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1976 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3952 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3951 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_494 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1976 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1975 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1974 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1973 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3953 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3954 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1977 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3954 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3953 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3955 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3956 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1978 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3956 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3955 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3957 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3958 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1979 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3958 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3957 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3959 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3960 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1980 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3960 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3959 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_495 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1980 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1979 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1978 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1977 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3961 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3962 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1981 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3962 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3961 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3963 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3964 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1982 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3964 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3963 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3965 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3966 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1983 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3966 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3965 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3967 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3968 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1984 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3968 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3967 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_496 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1984 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1983 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1982 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1981 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_124 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_496 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_495 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_494 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_493 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_31 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_124 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_123 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_122 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_121 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n8), .C(s83[1]), .D(n6), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n8), .C(s83[0]), .D(n6), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n7), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n7), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n7), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n7), .Z(sum8[0]) );
  CMX2X1 U3 ( .A0(n2), .A1(n3), .S(n6), .Z(n1) );
  CIVX2 U4 ( .A(n1), .Z(sum8[6]) );
  CMXI2X2 U5 ( .A0(n5), .A1(n4), .S(n8), .Z(sum8[7]) );
  CMX2X1 U6 ( .A0(c_out810), .A1(c_out811), .S(n8), .Z(c_out8) );
  CMXI2X1 U7 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n6) );
  CIVX2 U14 ( .A(n6), .Z(n8) );
  CIVX2 U15 ( .A(s83[2]), .Z(n3) );
  CIVX2 U16 ( .A(s84[2]), .Z(n2) );
  CIVX2 U17 ( .A(s83[3]), .Z(n5) );
  CIVX2 U18 ( .A(s84[3]), .Z(n4) );
  CIVX2 U19 ( .A(c_in8), .Z(n7) );
endmodule


module Add_half_3969 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3970 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1985 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3970 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3969 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3971 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3972 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1986 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3972 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3971 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3973 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3974 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1987 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3974 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3973 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3975 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3976 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1988 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3976 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3975 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_497 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1988 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1987 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1986 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1985 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3977 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3978 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1989 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3978 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3977 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3979 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3980 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1990 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3980 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3979 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3981 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3982 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1991 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3982 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3981 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3983 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3984 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1992 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3984 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3983 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_498 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1992 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1991 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1990 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1989 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3985 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3986 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1993 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3986 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3985 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3987 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3988 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1994 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3988 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3987 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3989 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3990 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1995 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3990 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3989 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3991 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3992 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_1996 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3992 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3991 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_499 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_1996 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1995 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1994 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1993 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_3993 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3994 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1997 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3994 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3993 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3995 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_3996 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1998 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3996 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3995 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3997 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_3998 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_1999 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_3998 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3997 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_3999 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4000 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2000 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4000 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_3999 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_500 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2000 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_1999 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_1998 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_1997 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_125 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_500 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_499 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_498 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_497 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_4001 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4002 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2001 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4002 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4001 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4003 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4004 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2002 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4004 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4003 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4005 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4006 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2003 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4006 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4005 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4007 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4008 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2004 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4008 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4007 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_501 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2004 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2003 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2002 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2001 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4009 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4010 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2005 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4010 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4009 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4011 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4012 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2006 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4012 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4011 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4013 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4014 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2007 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4014 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4013 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4015 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4016 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2008 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4016 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4015 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_502 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2008 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2007 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2006 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2005 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4017 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4018 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2009 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4018 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4017 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4019 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4020 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2010 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4020 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4019 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4021 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4022 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2011 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4022 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4021 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4023 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4024 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2012 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4024 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4023 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_503 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2012 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2011 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2010 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2009 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4025 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4026 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2013 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4026 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4025 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4027 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4028 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2014 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4028 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4027 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4029 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4030 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2015 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4030 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4029 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4031 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4032 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2016 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4032 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4031 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_504 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2016 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2015 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2014 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2013 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_126 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_504 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_503 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_502 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_501 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_4033 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4034 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2017 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4034 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4033 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4035 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4036 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2018 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4036 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4035 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4037 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4038 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2019 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4038 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4037 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4039 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4040 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2020 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4040 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4039 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_505 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2020 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2019 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2018 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2017 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4041 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4042 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2021 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4042 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4041 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4043 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4044 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2022 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4044 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4043 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4045 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4046 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2023 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4046 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4045 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4047 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4048 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2024 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4048 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4047 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_506 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2024 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2023 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2022 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2021 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4049 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4050 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2025 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4050 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4049 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4051 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4052 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2026 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4052 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4051 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4053 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4054 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2027 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4054 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4053 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4055 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4056 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2028 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4056 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4055 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_507 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2028 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2027 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2026 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2025 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4057 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4058 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2029 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4058 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4057 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4059 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4060 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2030 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4060 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4059 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4061 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4062 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2031 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4062 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4061 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4063 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4064 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2032 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4064 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4063 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_508 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2032 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2031 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2030 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2029 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_127 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_508 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_507 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_506 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_505 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_4065 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4066 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2033 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4066 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4065 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4067 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4068 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2034 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4068 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4067 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4069 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4070 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2035 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4070 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4069 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4071 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4072 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2036 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4072 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4071 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_509 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2036 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2035 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2034 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2033 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4073 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4074 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2037 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4074 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4073 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4075 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4076 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2038 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4076 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4075 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4077 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4078 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2039 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4078 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4077 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4079 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4080 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2040 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4080 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4079 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_510 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2040 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2039 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2038 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2037 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4081 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4082 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2041 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4082 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4081 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4083 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4084 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2042 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4084 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4083 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4085 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4086 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2043 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4086 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4085 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4087 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4088 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2044 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4088 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4087 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_511 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2044 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2043 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2042 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2041 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4089 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4090 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2045 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4090 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4089 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4091 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4092 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2046 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4092 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4091 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4093 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4094 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2047 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4094 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4093 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4095 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4096 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2048 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4096 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4095 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_512 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2048 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2047 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2046 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2045 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_128 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_512 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_511 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_510 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_509 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_32 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n4, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_128 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_127 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_126 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_125 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in8), .Z(n4) );
  CAOR2X1 U6 ( .A(s84[3]), .B(n5), .C(s83[3]), .D(n1), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n5), .C(s83[2]), .D(n1), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n5), .C(s83[1]), .D(n1), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n5), .C(s83[0]), .D(n1), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n4), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n4), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n4), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n4), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n5), .C(c_out810), .D(n1), .Z(c_out8) );
  CANR2X1 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n4), .Z(n1) );
endmodule


module bit32_8 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   c1, c2, c3;

  bit8_32 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8(a32[7:0]), .b8(b32[7:0]), 
        .c_in8(c_in32) );
  bit8_31 A322 ( .sum8(sum32[15:8]), .c_out8(c2), .a8(a32[15:8]), .b8(
        b32[15:8]), .c_in8(c1) );
  bit8_30 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8(a32[23:16]), .b8(
        b32[23:16]), .c_in8(c2) );
  bit8_29 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8(a32[31:24]), .b8(
        b32[31:24]), .c_in8(c3) );
endmodule


module Add_half_4097 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4098 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2049 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4098 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4097 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4099 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4100 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2050 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4100 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4099 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4101 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4102 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2051 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4102 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4101 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4103 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4104 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2052 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4104 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4103 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_513 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2052 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2051 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2050 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2049 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4105 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4106 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2053 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4106 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4105 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4107 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4108 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2054 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4108 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4107 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4109 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4110 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2055 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4110 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4109 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4111 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4112 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2056 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4112 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4111 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_514 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2056 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2055 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2054 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2053 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4113 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4114 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2057 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4114 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4113 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4115 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4116 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2058 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4116 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4115 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4117 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4118 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2059 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4118 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4117 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4119 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4120 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2060 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4120 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4119 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_515 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2060 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2059 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2058 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2057 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4121 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4122 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2061 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4122 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4121 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4123 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4124 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2062 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4124 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4123 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4125 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4126 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2063 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4126 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4125 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4127 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4128 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2064 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4128 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4127 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_516 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2064 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2063 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2062 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2061 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_129 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_516 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_515 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_514 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_513 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_4129 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4130 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2065 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4130 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4129 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4131 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4132 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2066 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4132 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4131 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4133 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4134 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2067 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4134 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4133 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4135 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4136 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2068 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4136 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4135 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_517 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2068 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2067 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2066 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2065 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4137 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4138 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2069 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4138 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4137 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4139 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4140 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2070 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4140 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4139 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4141 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4142 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2071 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4142 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4141 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4143 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4144 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2072 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4144 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4143 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_518 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2072 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2071 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2070 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2069 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4145 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4146 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2073 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4146 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4145 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4147 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4148 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2074 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4148 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4147 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4149 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4150 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2075 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4150 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4149 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4151 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4152 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2076 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4152 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4151 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_519 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2076 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2075 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2074 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2073 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4153 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4154 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2077 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4154 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4153 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4155 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4156 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2078 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4156 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4155 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4157 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4158 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2079 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4158 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4157 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4159 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4160 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2080 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4160 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4159 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_520 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2080 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2079 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2078 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2077 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_130 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_520 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_519 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_518 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_517 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_4161 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4162 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2081 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4162 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4161 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4163 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4164 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2082 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4164 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4163 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4165 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4166 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2083 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4166 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4165 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4167 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4168 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2084 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4168 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4167 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_521 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2084 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2083 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2082 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2081 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4169 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4170 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2085 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4170 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4169 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4171 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4172 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2086 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4172 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4171 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4173 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4174 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2087 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4174 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4173 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4175 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4176 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2088 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4176 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4175 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_522 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2088 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2087 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2086 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2085 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4177 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4178 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2089 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4178 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4177 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4179 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4180 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2090 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4180 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4179 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4181 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4182 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2091 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4182 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4181 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4183 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4184 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2092 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4184 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4183 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_523 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2092 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2091 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2090 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2089 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CAOR2XL U3 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CANR2X1 U6 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4185 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4186 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2093 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4186 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4185 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4187 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4188 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2094 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4188 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4187 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4189 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4190 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2095 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4190 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4189 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4191 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4192 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2096 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4192 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4191 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_524 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2096 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2095 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2094 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2093 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_131 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_524 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_523 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_522 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_521 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_4193 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4194 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2097 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4194 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4193 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4195 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4196 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2098 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4196 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4195 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4197 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4198 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2099 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4198 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4197 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4199 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4200 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2100 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4200 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4199 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_525 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2100 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2099 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2098 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2097 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CAOR2XL U3 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CANR2X1 U6 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4201 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4202 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2101 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4202 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4201 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4203 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4204 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2102 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4204 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4203 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4205 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4206 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2103 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4206 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4205 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4207 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4208 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2104 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4208 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4207 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_526 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2104 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2103 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2102 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2101 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4209 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4210 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2105 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4210 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4209 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4211 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4212 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2106 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4212 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4211 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4213 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4214 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2107 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4214 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4213 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4215 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4216 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2108 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4216 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4215 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_527 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2108 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2107 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2106 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2105 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CAOR2XL U3 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CANR2X1 U6 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4217 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4218 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2109 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4218 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4217 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4219 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4220 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2110 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4220 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4219 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4221 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4222 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2111 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4222 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4221 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4223 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4224 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2112 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4224 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4223 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_528 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2112 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2111 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2110 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2109 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_132 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_528 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_527 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_526 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_525 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_33 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n3, n4, n5, n6;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_132 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_131 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_130 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_129 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X2 U3 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2X2 U4 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2X2 U5 ( .A0(s83[0]), .A1(s84[0]), .S(n6), .Z(sum8[4]) );
  CMX2X1 U6 ( .A0(s83[3]), .A1(s84[3]), .S(n6), .Z(sum8[7]) );
  CMX2X1 U7 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2X2 U8 ( .A0(s81[0]), .A1(s82[0]), .S(c_in8), .Z(sum8[0]) );
  CMX2X1 U9 ( .A0(s83[2]), .A1(s84[2]), .S(n6), .Z(sum8[6]) );
  CMX2X1 U10 ( .A0(s83[1]), .A1(s84[1]), .S(n6), .Z(sum8[5]) );
  CIVX2 U11 ( .A(n3), .Z(n6) );
  CIVX2 U12 ( .A(c_out810), .Z(n5) );
  CIVX2 U13 ( .A(c_out811), .Z(n4) );
  CMXI2X1 U14 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n3) );
  CMXI2X1 U15 ( .A0(n5), .A1(n4), .S(n6), .Z(c_out8) );
endmodule


module Add_half_4225 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4226 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2113 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4226 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4225 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4227 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4228 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2114 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4228 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4227 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4229 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4230 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2115 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4230 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4229 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4231 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4232 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2116 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4232 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4231 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_529 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2116 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2115 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2114 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2113 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_4233 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4234 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2117 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4234 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4233 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4235 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4236 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2118 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4236 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4235 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4237 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4238 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2119 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4238 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4237 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4239 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4240 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2120 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4240 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4239 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_530 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2120 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2119 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2118 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2117 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CIVXL U3 ( .A(s3), .Z(n4) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_4241 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4242 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2121 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4242 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4241 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4243 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4244 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2122 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4244 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4243 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4245 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4246 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2123 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4246 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4245 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4247 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4248 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2124 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4248 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4247 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_531 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2124 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2123 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2122 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2121 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_4249 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4250 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2125 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4250 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4249 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4251 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4252 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2126 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4252 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4251 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4253 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4254 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2127 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4254 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4253 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4255 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4256 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2128 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4256 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4255 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_532 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2128 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2127 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2126 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2125 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVXL U3 ( .A(s3), .Z(n6) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module bit4_133 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_532 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_531 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_530 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_529 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n3), .Z(sum4[0]) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n2), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n2), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(c_out410), .A1(c_out411), .S(n2), .Z(c_out4) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMXI2X1 U7 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n2) );
  CIVX2 U10 ( .A(c_in4), .Z(n3) );
endmodule


module Add_half_4257 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4258 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2129 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4258 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4257 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4259 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4260 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2130 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4260 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4259 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4261 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4262 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2131 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4262 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4261 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4263 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4264 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2132 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4264 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4263 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_533 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2132 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2131 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2130 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2129 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_4265 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4266 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2133 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4266 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4265 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4267 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4268 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2134 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4268 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4267 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4269 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4270 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2135 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4270 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4269 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4271 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4272 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2136 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4272 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4271 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_534 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2136 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2135 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2134 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2133 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4273 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4274 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2137 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4274 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4273 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4275 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4276 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2138 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4276 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4275 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4277 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4278 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2139 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4278 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4277 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4279 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4280 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2140 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4280 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4279 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_535 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2140 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2139 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2138 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2137 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_4281 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4282 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2141 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4282 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4281 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4283 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4284 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2142 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4284 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4283 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4285 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4286 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2143 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4286 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4285 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4287 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4288 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2144 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4288 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4287 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_536 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2144 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2143 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2142 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2141 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module bit4_134 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_536 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_535 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_534 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_533 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n11), .Z(sum4[0]) );
  CIVX2 U3 ( .A(c_out410), .Z(n3) );
  CIVX2 U4 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n8) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U8 ( .A(s41[1]), .Z(n5) );
  CIVX2 U10 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(s43[0]), .Z(n7) );
  CIVX2 U13 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX2 U15 ( .A(s43[1]), .Z(n10) );
  CIVX2 U16 ( .A(s44[1]), .Z(n9) );
  CMXI2X1 U17 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
  CIVX2 U18 ( .A(c_in4), .Z(n11) );
endmodule


module Add_half_4289 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4290 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2145 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4290 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4289 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4291 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4292 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2146 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4292 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4291 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4293 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4294 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2147 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4294 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4293 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4295 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4296 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2148 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4296 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4295 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_537 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2148 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2147 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2146 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2145 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(n1), .Z(n2) );
  CIVX2 U6 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_4297 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4298 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2149 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4298 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4297 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4299 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4300 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2150 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4300 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4299 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4301 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4302 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2151 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4302 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4301 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4303 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4304 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2152 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4304 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4303 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_538 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2152 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2151 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2150 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2149 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CIVXL U3 ( .A(s3), .Z(n4) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_4305 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4306 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2153 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4306 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4305 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4307 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4308 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2154 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4308 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4307 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4309 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4310 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2155 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4310 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4309 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4311 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4312 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2156 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4312 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4311 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_539 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2156 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2155 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2154 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2153 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_4313 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4314 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2157 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4314 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4313 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4315 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4316 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2158 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4316 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4315 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4317 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4318 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2159 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4318 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4317 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4319 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4320 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2160 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4320 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4319 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_540 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2160 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2159 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2158 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2157 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(s3), .Z(n6) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module bit4_135 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_540 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_539 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_538 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_537 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n6), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n6), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n6) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out4) );
  CIVX2 U11 ( .A(s41[0]), .Z(n5) );
  CIVX2 U12 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
endmodule


module Add_half_4321 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4322 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2161 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4322 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4321 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4323 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4324 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2162 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4324 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4323 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4325 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4326 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2163 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4326 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4325 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4327 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4328 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2164 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4328 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4327 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_541 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_2164 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2163 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2162 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2161 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_4329 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4330 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2165 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4330 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4329 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4331 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4332 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2166 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4332 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4331 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4333 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4334 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2167 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4334 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4333 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4335 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4336 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2168 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4336 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4335 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_542 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_2168 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2167 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2166 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2165 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_4337 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4338 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2169 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4338 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4337 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4339 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4340 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2170 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4340 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4339 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4341 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4342 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2171 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4342 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4341 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4343 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4344 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2172 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4344 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4343 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_543 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2172 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2171 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2170 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2169 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_4345 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4346 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2173 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4346 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4345 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4347 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4348 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2174 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4348 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4347 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4349 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_4350 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2175 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4350 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4349 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4351 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4352 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2176 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4352 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4351 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_544 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2176 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2175 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2174 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2173 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_136 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_544 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_543 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_542 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_541 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U4 ( .A(c_out410), .Z(n3) );
  CIVX2 U5 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n8) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U9 ( .A(s41[1]), .Z(n5) );
  CIVX2 U10 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(s43[0]), .Z(n7) );
  CIVX2 U13 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX2 U15 ( .A(s43[1]), .Z(n10) );
  CIVX2 U16 ( .A(s44[1]), .Z(n9) );
  CMXI2X1 U17 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
endmodule


module bit8_34 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_136 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_135 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_134 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_133 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVXL U3 ( .A(c_in8), .Z(n1) );
  CIVXL U4 ( .A(n1), .Z(n2) );
  CMX2X1 U5 ( .A0(s83[0]), .A1(s84[0]), .S(n3), .Z(sum8[4]) );
  CMX2X2 U6 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n3) );
  CMX2X1 U7 ( .A0(s81[0]), .A1(s82[0]), .S(c_in8), .Z(sum8[0]) );
  CMX2X2 U8 ( .A0(c_out810), .A1(c_out811), .S(n3), .Z(c_out8) );
  CMX2X1 U9 ( .A0(s83[2]), .A1(s84[2]), .S(n3), .Z(sum8[6]) );
  CMX2X1 U10 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2X1 U11 ( .A0(s81[3]), .A1(s82[3]), .S(n2), .Z(sum8[3]) );
  CMX2X1 U12 ( .A0(s83[3]), .A1(s84[3]), .S(n3), .Z(sum8[7]) );
  CMX2X1 U13 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2X1 U14 ( .A0(s83[1]), .A1(s84[1]), .S(n3), .Z(sum8[5]) );
endmodule


module Add_half_4353 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4354 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2177 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4354 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4353 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4355 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4356 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2178 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4356 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4355 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4357 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4358 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2179 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4358 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4357 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4359 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4360 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2180 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4360 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4359 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_545 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2180 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2179 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2178 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2177 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(s4), .Z(n5) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CIVX2 U7 ( .A(s1), .Z(n3) );
  CIVX2 U8 ( .A(s2), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_4361 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4362 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2181 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4362 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4361 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4363 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4364 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2182 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4364 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4363 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4365 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_4366 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2183 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4366 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4365 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4367 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4368 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2184 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4368 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4367 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_546 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2184 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2183 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2182 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2181 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_4369 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4370 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENXL U1 ( .A(a), .B(b), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2185 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4370 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4369 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4371 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4372 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2186 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4372 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4371 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4373 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4374 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2187 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_4374 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4373 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_4375 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4376 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2188 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4376 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4375 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_547 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_2188 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2187 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2186 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2185 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(c_out10), .Z(n3) );
  CIVX1 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_4377 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(a), .B(n2), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_4378 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2189 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4378 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4377 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4379 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4380 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX1 U1 ( .A(a), .B(b), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2190 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4380 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4379 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4381 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_4382 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2191 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_4382 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4381 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_4383 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4384 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2192 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_4384 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4383 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_548 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2192 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2191 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2190 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2189 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX1 U4 ( .A(n1), .Z(n4) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2XL U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_137 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_548 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_547 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_546 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_545 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n2) );
  CMX2XL U4 ( .A0(s43[1]), .A1(s44[1]), .S(n2), .Z(sum4[3]) );
  CMX2XL U5 ( .A0(s43[0]), .A1(s44[0]), .S(n2), .Z(sum4[2]) );
  CMX2X1 U6 ( .A0(c_out410), .A1(c_out411), .S(n2), .Z(c_out4) );
  CMX2X1 U7 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U8 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
endmodule


module Add_half_4385 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4386 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2193 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4386 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4385 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4387 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4388 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2194 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4388 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4387 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4389 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4390 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2195 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4390 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4389 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4391 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4392 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2196 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4392 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4391 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_549 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_2196 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2195 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2194 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2193 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_4393 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4394 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2197 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4394 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4393 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4395 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4396 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2198 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4396 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4395 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4397 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4398 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2199 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_4398 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4397 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4399 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4400 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2200 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_4400 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4399 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X2 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_550 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_2200 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2199 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2198 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2197 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2X1 U4 ( .A0(c_out11), .A1(c_out10), .S(n2), .Z(c_out2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module Add_half_4401 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4402 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2201 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4402 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4401 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4403 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4404 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2202 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4404 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4403 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4405 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4406 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2203 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4406 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4405 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4407 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4408 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2204 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_4408 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4407 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CND2X1 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_551 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_2204 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2203 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2202 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2201 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
endmodule


module Add_half_4409 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4410 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2205 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4410 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4409 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4411 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4412 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2206 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4412 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4411 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4413 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4414 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2207 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_4414 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4413 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CND2X1 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_4415 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4416 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2208 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_4416 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4415 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CND2X1 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_552 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2208 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2207 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2206 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2205 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(c_out11), .Z(n2) );
  CIVX1 U4 ( .A(c_out10), .Z(n3) );
  CIVX1 U5 ( .A(n1), .Z(n4) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_138 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_552 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_551 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_550 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_549 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVXL U3 ( .A(n2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CIVXL U5 ( .A(s42[1]), .Z(n7) );
  CMXI2XL U6 ( .A0(n13), .A1(n12), .S(n1), .Z(sum4[3]) );
  CIVX1 U7 ( .A(s42[0]), .Z(n5) );
  CIVX1 U8 ( .A(s41[0]), .Z(n6) );
  CIVX2 U9 ( .A(c_out410), .Z(n4) );
  CIVX2 U10 ( .A(c_out411), .Z(n3) );
  CIVX2 U11 ( .A(n2), .Z(n11) );
  CMXI2X1 U12 ( .A0(n4), .A1(n3), .S(n11), .Z(c_out4) );
  CMXI2X1 U13 ( .A0(n6), .A1(n5), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U14 ( .A(s41[1]), .Z(n8) );
  CMXI2X1 U15 ( .A0(n8), .A1(n7), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U16 ( .A(s43[0]), .Z(n10) );
  CIVX2 U17 ( .A(s44[0]), .Z(n9) );
  CMXI2X1 U18 ( .A0(n10), .A1(n9), .S(n11), .Z(sum4[2]) );
  CIVX2 U19 ( .A(s43[1]), .Z(n13) );
  CIVX2 U20 ( .A(s44[1]), .Z(n12) );
endmodule


module Add_half_4417 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4418 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2209 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4418 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4417 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4419 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4420 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2210 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4420 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4419 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4421 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4422 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2211 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4422 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4421 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4423 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4424 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2212 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4424 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4423 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_553 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2212 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2211 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2210 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2209 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4425 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4426 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2213 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4426 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4425 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4427 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4428 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2214 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4428 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4427 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4429 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4430 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2215 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4430 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4429 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4431 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4432 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2216 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4432 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4431 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_554 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2216 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2215 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2214 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2213 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4433 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4434 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2217 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4434 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4433 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4435 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4436 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2218 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4436 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4435 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4437 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4438 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2219 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4438 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4437 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4439 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4440 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2220 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4440 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4439 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_555 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2220 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2219 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2218 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2217 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4441 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4442 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2221 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4442 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4441 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4443 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4444 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2222 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4444 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4443 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4445 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4446 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2223 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4446 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4445 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4447 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4448 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2224 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4448 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4447 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_556 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2224 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2223 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2222 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2221 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_139 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_556 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_555 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_554 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_553 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_4449 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4450 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2225 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4450 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4449 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4451 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4452 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2226 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4452 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4451 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4453 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4454 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2227 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4454 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4453 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4455 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4456 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2228 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4456 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4455 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_557 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2228 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2227 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2226 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2225 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4457 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4458 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2229 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4458 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4457 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4459 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4460 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2230 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4460 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4459 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4461 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4462 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2231 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4462 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4461 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4463 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4464 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2232 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4464 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4463 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_558 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2232 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2231 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2230 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2229 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4465 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4466 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2233 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4466 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4465 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4467 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4468 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2234 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4468 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4467 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4469 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4470 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2235 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4470 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4469 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4471 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4472 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2236 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4472 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4471 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_559 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2236 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2235 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2234 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2233 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4473 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4474 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2237 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4474 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4473 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4475 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4476 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2238 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4476 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4475 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4477 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4478 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2239 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4478 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4477 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4479 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4480 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2240 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4480 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4479 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_560 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2240 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2239 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2238 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2237 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_140 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_560 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_559 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_558 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_557 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_35 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_140 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_139 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_138 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_137 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n7), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n7), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n7), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n7), .Z(sum8[0]) );
  CMXI2X2 U3 ( .A0(n3), .A1(n2), .S(n6), .Z(sum8[4]) );
  CMXI2X2 U4 ( .A0(n5), .A1(n4), .S(n6), .Z(sum8[5]) );
  CMX2X2 U5 ( .A0(c_out811), .A1(c_out810), .S(n1), .Z(c_out8) );
  CIVX1 U6 ( .A(s83[1]), .Z(n5) );
  CMX2X2 U7 ( .A0(s83[2]), .A1(s84[2]), .S(n6), .Z(sum8[6]) );
  CMX2X2 U8 ( .A0(s83[3]), .A1(s84[3]), .S(n6), .Z(sum8[7]) );
  CMXI2X1 U9 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CIVX2 U14 ( .A(n1), .Z(n6) );
  CIVX2 U15 ( .A(s83[0]), .Z(n3) );
  CIVX2 U16 ( .A(s84[0]), .Z(n2) );
  CIVX2 U17 ( .A(s84[1]), .Z(n4) );
  CIVX2 U18 ( .A(c_in8), .Z(n7) );
endmodule


module Add_half_4481 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4482 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2241 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4482 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4481 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4483 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4484 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2242 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4484 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4483 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4485 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4486 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2243 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4486 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4485 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4487 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4488 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2244 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4488 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4487 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_561 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2244 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2243 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2242 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2241 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4489 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4490 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2245 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4490 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4489 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4491 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4492 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2246 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4492 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4491 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4493 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4494 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2247 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4494 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4493 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4495 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4496 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2248 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4496 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4495 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_562 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2248 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2247 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2246 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2245 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4497 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4498 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2249 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4498 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4497 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4499 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4500 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2250 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4500 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4499 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4501 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4502 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2251 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4502 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4501 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4503 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4504 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2252 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4504 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4503 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_563 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2252 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2251 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2250 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2249 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4505 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4506 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2253 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4506 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4505 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4507 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4508 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2254 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4508 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4507 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4509 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4510 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2255 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4510 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4509 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4511 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4512 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2256 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4512 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4511 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_564 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2256 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2255 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2254 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2253 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_141 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_564 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_563 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_562 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_561 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_4513 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4514 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2257 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4514 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4513 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4515 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4516 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2258 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4516 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4515 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4517 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4518 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2259 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4518 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4517 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4519 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4520 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2260 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4520 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4519 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_565 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2260 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2259 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2258 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2257 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4521 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4522 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2261 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4522 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4521 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4523 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4524 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2262 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4524 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4523 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4525 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4526 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2263 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4526 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4525 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4527 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4528 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2264 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4528 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4527 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_566 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2264 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2263 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2262 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2261 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4529 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4530 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2265 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4530 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4529 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4531 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4532 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2266 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4532 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4531 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4533 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4534 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2267 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4534 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4533 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4535 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4536 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2268 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4536 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4535 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_567 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2268 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2267 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2266 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2265 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4537 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4538 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2269 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4538 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4537 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4539 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4540 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2270 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4540 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4539 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4541 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4542 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2271 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4542 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4541 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4543 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4544 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2272 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4544 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4543 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_568 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2272 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2271 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2270 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2269 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_142 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_568 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_567 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_566 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_565 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_4545 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4546 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2273 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4546 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4545 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4547 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4548 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2274 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4548 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4547 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4549 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4550 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2275 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4550 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4549 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4551 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4552 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2276 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4552 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4551 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_569 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2276 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2275 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2274 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2273 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4553 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4554 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2277 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4554 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4553 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4555 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4556 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2278 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4556 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4555 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4557 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4558 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2279 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4558 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4557 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4559 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4560 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2280 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4560 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4559 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_570 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2280 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2279 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2278 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2277 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4561 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4562 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2281 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4562 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4561 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4563 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4564 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2282 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4564 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4563 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4565 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4566 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2283 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4566 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4565 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4567 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4568 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2284 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4568 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4567 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_571 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2284 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2283 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2282 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2281 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4569 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4570 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2285 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4570 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4569 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4571 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4572 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2286 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4572 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4571 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4573 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4574 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2287 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4574 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4573 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4575 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4576 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2288 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4576 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4575 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_572 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2288 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2287 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2286 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2285 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_143 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_572 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_571 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_570 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_569 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_4577 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4578 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2289 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4578 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4577 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4579 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4580 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2290 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4580 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4579 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4581 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4582 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2291 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4582 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4581 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4583 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4584 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2292 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4584 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4583 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_573 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2292 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2291 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2290 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2289 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4585 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4586 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2293 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4586 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4585 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4587 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4588 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2294 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4588 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4587 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4589 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4590 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2295 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4590 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4589 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4591 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4592 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2296 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4592 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4591 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_574 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2296 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2295 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2294 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2293 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4593 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4594 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2297 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4594 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4593 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4595 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4596 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2298 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4596 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4595 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4597 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4598 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2299 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4598 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4597 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4599 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4600 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2300 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4600 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4599 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_575 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2300 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2299 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2298 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2297 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4601 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4602 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2301 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4602 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4601 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4603 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4604 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2302 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4604 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4603 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4605 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4606 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2303 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4606 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4605 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4607 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4608 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2304 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4608 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4607 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_576 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2304 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2303 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2302 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2301 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_144 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_576 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_575 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_574 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_573 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_36 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n4, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_144 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_143 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_142 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_141 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in8), .Z(n4) );
  CAOR2X1 U6 ( .A(s84[3]), .B(n5), .C(s83[3]), .D(n1), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n5), .C(s83[2]), .D(n1), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n5), .C(s83[1]), .D(n1), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n5), .C(s83[0]), .D(n1), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n4), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n4), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n4), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n4), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n5), .C(c_out810), .D(n1), .Z(c_out8) );
  CANR2X1 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n4), .Z(n1) );
endmodule


module bit32_9 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   c1, c2, c3;

  bit8_36 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8(a32[7:0]), .b8(b32[7:0]), 
        .c_in8(c_in32) );
  bit8_35 A322 ( .sum8(sum32[15:8]), .c_out8(c2), .a8(a32[15:8]), .b8(
        b32[15:8]), .c_in8(c1) );
  bit8_34 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8(a32[23:16]), .b8(
        b32[23:16]), .c_in8(c2) );
  bit8_33 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8(a32[31:24]), .b8(
        b32[31:24]), .c_in8(c3) );
endmodule


module Add_half_4609 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4610 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2305 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4610 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4609 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4611 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4612 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2306 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4612 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4611 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4613 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4614 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2307 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4614 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4613 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4615 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4616 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2308 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4616 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4615 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_577 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2308 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2307 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2306 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2305 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4617 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4618 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2309 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4618 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4617 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4619 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4620 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2310 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4620 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4619 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4621 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4622 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2311 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4622 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4621 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4623 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4624 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2312 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4624 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4623 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_578 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2312 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2311 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2310 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2309 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4625 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4626 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2313 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4626 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4625 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4627 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4628 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2314 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4628 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4627 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4629 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4630 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2315 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4630 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4629 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4631 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4632 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2316 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4632 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4631 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_579 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2316 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2315 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2314 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2313 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4633 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4634 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2317 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4634 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4633 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4635 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4636 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2318 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4636 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4635 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4637 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4638 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2319 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4638 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4637 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4639 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4640 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2320 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4640 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4639 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_580 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2320 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2319 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2318 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2317 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_145 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_580 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_579 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_578 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_577 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_4641 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4642 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2321 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4642 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4641 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4643 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4644 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2322 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4644 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4643 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4645 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4646 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2323 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4646 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4645 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4647 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4648 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2324 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4648 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4647 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_581 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2324 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2323 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2322 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2321 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4649 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4650 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2325 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4650 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4649 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4651 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4652 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2326 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4652 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4651 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4653 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4654 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2327 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4654 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4653 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4655 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4656 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2328 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4656 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4655 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_582 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2328 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2327 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2326 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2325 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4657 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4658 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2329 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4658 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4657 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4659 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4660 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2330 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4660 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4659 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4661 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4662 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2331 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4662 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4661 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4663 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4664 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2332 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4664 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4663 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_583 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2332 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2331 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2330 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2329 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4665 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4666 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2333 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4666 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4665 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4667 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4668 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2334 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4668 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4667 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4669 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4670 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2335 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4670 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4669 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4671 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4672 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2336 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4672 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4671 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_584 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2336 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2335 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2334 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2333 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_146 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_584 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_583 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_582 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_581 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_4673 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4674 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2337 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4674 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4673 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4675 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4676 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2338 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4676 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4675 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4677 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4678 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2339 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4678 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4677 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4679 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4680 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2340 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4680 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4679 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_585 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2340 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2339 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2338 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2337 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4681 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4682 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2341 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4682 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4681 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4683 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4684 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2342 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4684 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4683 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4685 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4686 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2343 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4686 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4685 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4687 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4688 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2344 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4688 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4687 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_586 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2344 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2343 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2342 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2341 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4689 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4690 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2345 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4690 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4689 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4691 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4692 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2346 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4692 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4691 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4693 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4694 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2347 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4694 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4693 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4695 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4696 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2348 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4696 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4695 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_587 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2348 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2347 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2346 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2345 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CAOR2XL U3 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CANR2X1 U7 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4697 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4698 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2349 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4698 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4697 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4699 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4700 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2350 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4700 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4699 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4701 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4702 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2351 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4702 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4701 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4703 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4704 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2352 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4704 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4703 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_588 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2352 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2351 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2350 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2349 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_147 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_588 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_587 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_586 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_585 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
endmodule


module Add_half_4705 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4706 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2353 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4706 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4705 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4707 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4708 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2354 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4708 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4707 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4709 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4710 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2355 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4710 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4709 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4711 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4712 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2356 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4712 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4711 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_589 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2356 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2355 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2354 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2353 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CAOR2XL U3 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2XL U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CANR2X1 U7 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4713 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4714 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2357 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4714 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4713 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4715 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4716 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2358 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4716 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4715 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4717 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4718 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2359 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4718 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4717 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4719 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4720 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2360 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4720 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4719 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_590 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2360 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2359 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2358 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2357 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4721 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4722 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2361 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4722 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4721 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4723 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4724 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2362 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4724 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4723 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4725 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4726 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2363 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4726 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4725 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4727 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4728 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2364 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4728 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4727 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_591 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2364 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2363 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2362 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2361 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CAOR2XL U3 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CANR2X1 U6 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4729 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4730 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2365 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4730 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4729 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4731 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4732 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2366 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4732 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4731 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4733 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4734 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2367 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4734 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4733 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4735 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4736 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2368 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4736 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4735 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_592 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2368 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2367 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2366 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2365 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_148 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_592 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_591 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_590 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_589 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2XL U3 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X2 U10 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_37 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_148 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_147 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_146 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_145 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X4 U3 ( .A0(s81[0]), .A1(s82[0]), .S(c_in8), .Z(sum8[0]) );
  CMXI2XL U4 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out8) );
  CMX2X2 U5 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2X4 U6 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2X2 U7 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CMX2X2 U8 ( .A0(s83[0]), .A1(s84[0]), .S(n1), .Z(sum8[4]) );
  CMX2XL U9 ( .A0(s83[3]), .A1(s84[3]), .S(n1), .Z(sum8[7]) );
  CMX2X1 U10 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2X1 U11 ( .A0(s83[2]), .A1(s84[2]), .S(n1), .Z(sum8[6]) );
  CMX2X1 U12 ( .A0(s83[1]), .A1(s84[1]), .S(n1), .Z(sum8[5]) );
  CIVX2 U13 ( .A(c_out810), .Z(n3) );
  CIVX2 U14 ( .A(c_out811), .Z(n2) );
endmodule


module Add_half_4737 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4738 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2369 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4738 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4737 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4739 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4740 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2370 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4740 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4739 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4741 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4742 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2371 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4742 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4741 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4743 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4744 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2372 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4744 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4743 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_593 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2372 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2371 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2370 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2369 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_4745 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4746 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2373 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4746 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4745 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4747 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4748 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2374 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4748 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4747 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4749 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4750 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2375 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4750 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4749 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4751 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4752 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2376 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4752 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4751 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_594 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2376 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2375 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2374 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2373 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CIVXL U3 ( .A(s3), .Z(n4) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_4753 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4754 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2377 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4754 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4753 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4755 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4756 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2378 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4756 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4755 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4757 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4758 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2379 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4758 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4757 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4759 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4760 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2380 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4760 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4759 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_595 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2380 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2379 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2378 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2377 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_4761 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4762 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2381 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4762 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4761 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4763 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4764 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2382 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4764 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4763 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4765 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4766 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2383 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4766 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4765 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4767 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4768 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2384 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4768 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4767 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_596 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2384 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2383 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2382 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2381 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX1 U3 ( .A(s3), .Z(n6) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module bit4_149 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_596 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_595 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_594 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_593 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n5), .Z(sum4[0]) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2X1 U4 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
  CIVX2 U12 ( .A(c_in4), .Z(n5) );
endmodule


module Add_half_4769 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4770 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2385 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4770 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4769 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4771 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4772 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2386 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4772 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4771 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4773 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4774 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2387 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4774 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4773 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4775 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4776 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2388 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4776 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4775 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_597 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2388 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2387 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2386 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2385 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_4777 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4778 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2389 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4778 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4777 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4779 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4780 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2390 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4780 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4779 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4781 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4782 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2391 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4782 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4781 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4783 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4784 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2392 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4784 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4783 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_598 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2392 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2391 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2390 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2389 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4785 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4786 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2393 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4786 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4785 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4787 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4788 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2394 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4788 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4787 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4789 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4790 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2395 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4790 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4789 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4791 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4792 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2396 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4792 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4791 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_599 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2396 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2395 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2394 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2393 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_4793 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4794 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2397 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4794 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4793 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4795 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4796 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2398 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4796 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4795 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4797 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4798 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2399 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4798 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4797 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4799 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4800 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2400 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4800 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4799 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_600 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2400 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2399 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2398 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2397 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module bit4_150 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_600 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_599 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_598 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_597 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n11), .Z(sum4[0]) );
  CIVX2 U3 ( .A(c_out410), .Z(n3) );
  CIVX2 U4 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n8) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U8 ( .A(s41[1]), .Z(n5) );
  CIVX2 U10 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(s43[0]), .Z(n7) );
  CIVX2 U13 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX2 U15 ( .A(s43[1]), .Z(n10) );
  CIVX2 U16 ( .A(s44[1]), .Z(n9) );
  CMXI2X1 U17 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
  CIVX2 U18 ( .A(c_in4), .Z(n11) );
endmodule


module Add_half_4801 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4802 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2401 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4802 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4801 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4803 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4804 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2402 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4804 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4803 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4805 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4806 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2403 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4806 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4805 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4807 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4808 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2404 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4808 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4807 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_601 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2404 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2403 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2402 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2401 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(n1), .Z(n2) );
  CIVX2 U6 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_4809 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4810 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2405 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4810 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4809 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4811 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4812 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2406 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4812 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4811 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4813 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4814 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2407 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4814 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4813 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4815 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4816 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2408 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4816 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4815 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_602 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2408 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2407 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2406 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2405 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CIVX1 U3 ( .A(s3), .Z(n4) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_4817 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4818 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2409 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4818 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4817 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4819 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4820 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2410 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4820 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4819 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4821 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4822 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2411 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4822 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4821 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4823 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4824 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2412 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4824 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4823 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_603 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_2412 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2411 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2410 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2409 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_4825 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4826 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2413 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4826 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4825 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4827 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4828 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2414 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4828 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4827 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4829 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_4830 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2415 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4830 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4829 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4831 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4832 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2416 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4832 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4831 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_604 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2416 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2415 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2414 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2413 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(s3), .Z(n6) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module bit4_151 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_604 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_603 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_602 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_601 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module Add_half_4833 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4834 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2417 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4834 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4833 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4835 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4836 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2418 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4836 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4835 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4837 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4838 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2419 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4838 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4837 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4839 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4840 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2420 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4840 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4839 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_605 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_2420 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2419 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2418 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2417 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_4841 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4842 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2421 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4842 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4841 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4843 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4844 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2422 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4844 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4843 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4845 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4846 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2423 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4846 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4845 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4847 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4848 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2424 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4848 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4847 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_606 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_2424 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2423 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2422 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2421 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_4849 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4850 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2425 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4850 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4849 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4851 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4852 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2426 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4852 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4851 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4853 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4854 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2427 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4854 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4853 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4855 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4856 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2428 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4856 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4855 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_607 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2428 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2427 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2426 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2425 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_4857 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4858 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2429 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4858 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4857 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4859 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4860 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2430 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4860 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4859 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4861 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4862 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2431 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4862 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4861 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4863 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4864 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2432 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4864 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4863 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_608 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2432 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2431 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2430 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2429 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_152 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_608 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_607 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_606 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_605 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(c_out410), .Z(n3) );
  CIVX2 U4 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n10) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n10), .Z(c_out4) );
  CIVX2 U8 ( .A(s41[0]), .Z(n5) );
  CIVX2 U9 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U11 ( .A(s41[1]), .Z(n7) );
  CIVX2 U12 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U13 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n9) );
  CIVX2 U15 ( .A(s44[0]), .Z(n8) );
  CMXI2X1 U16 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CIVX2 U17 ( .A(s43[1]), .Z(n12) );
  CIVX2 U18 ( .A(s44[1]), .Z(n11) );
  CMXI2X1 U19 ( .A0(n12), .A1(n11), .S(n10), .Z(sum4[3]) );
endmodule


module bit8_38 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_152 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_151 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_150 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_149 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2XL U3 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2X2 U4 ( .A0(c_out810), .A1(c_out811), .S(n8), .Z(c_out8) );
  CIVX2 U5 ( .A(n1), .Z(n8) );
  CMXI2X1 U6 ( .A0(n5), .A1(n4), .S(n8), .Z(sum8[4]) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(c_in8), .Z(sum8[0]) );
  CMX2X1 U8 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2X1 U9 ( .A0(s83[3]), .A1(s84[3]), .S(n8), .Z(sum8[7]) );
  CMX2X1 U10 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2X1 U11 ( .A0(s83[1]), .A1(s84[1]), .S(n8), .Z(sum8[5]) );
  CMXI2X2 U12 ( .A0(n7), .A1(n6), .S(n8), .Z(sum8[6]) );
  CMXI2X1 U13 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CIVX2 U14 ( .A(s81[0]), .Z(n3) );
  CIVX2 U15 ( .A(s82[0]), .Z(n2) );
  CIVX2 U16 ( .A(s83[0]), .Z(n5) );
  CIVX2 U17 ( .A(s84[0]), .Z(n4) );
  CIVX2 U18 ( .A(s83[2]), .Z(n7) );
  CIVX2 U19 ( .A(s84[2]), .Z(n6) );
endmodule


module Add_half_4865 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_4866 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2433 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4866 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4865 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4867 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4868 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2434 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4868 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4867 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4869 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_4870 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2435 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4870 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4869 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4871 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4872 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2436 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4872 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4871 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_609 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_2436 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2435 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2434 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2433 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_4873 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4874 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2437 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4874 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4873 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4875 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4876 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2438 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4876 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4875 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4877 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4878 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2439 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4878 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4877 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4879 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4880 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2440 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4880 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4879 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_610 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2440 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2439 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2438 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2437 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(n1), .Z(n4) );
  CIVX2 U6 ( .A(s1), .Z(n3) );
  CIVX2 U7 ( .A(s2), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_4881 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4882 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2441 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4882 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4881 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4883 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4884 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2442 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4884 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4883 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4885 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4886 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2443 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4886 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4885 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4887 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4888 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2444 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4888 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4887 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_611 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2444 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2443 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2442 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2441 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_4889 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4890 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2445 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4890 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4889 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4891 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4892 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2446 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4892 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4891 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4893 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4894 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2447 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4894 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4893 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4895 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4896 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2448 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4896 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4895 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_612 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2448 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2447 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2446 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2445 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_153 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_612 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_611 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_610 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_609 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n8), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n8), .Z(sum4[2]) );
  CIVX1 U5 ( .A(c_out410), .Z(n3) );
  CIVX2 U6 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n8) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U10 ( .A(s41[0]), .Z(n5) );
  CIVX2 U11 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U13 ( .A(s41[1]), .Z(n7) );
  CIVX2 U14 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U15 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
endmodule


module Add_half_4897 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4898 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2449 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4898 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4897 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4899 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4900 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2450 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4900 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4899 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4901 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4902 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2451 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4902 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4901 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4903 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4904 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2452 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4904 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4903 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_613 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2452 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2451 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2450 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2449 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_4905 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4906 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2453 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4906 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4905 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4907 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4908 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2454 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4908 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4907 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4909 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4910 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2455 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4910 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4909 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4911 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4912 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2456 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4912 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4911 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_614 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_2456 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2455 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2454 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2453 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_4913 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_4914 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2457 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4914 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4913 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4915 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4916 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2458 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4916 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4915 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4917 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4918 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2459 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4918 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4917 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4919 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4920 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2460 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_4920 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4919 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_615 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2460 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2459 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2458 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2457 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s1), .Z(n5) );
  CMXI2X1 U4 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n6) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_4921 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4922 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2461 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4922 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4921 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4923 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4924 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2462 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4924 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4923 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4925 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_4926 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2463 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_4926 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4925 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4927 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4928 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2464 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4928 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4927 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_616 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2464 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2463 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2462 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2461 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module bit4_154 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_616 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_615 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_614 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_613 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n6), .A1(n5), .S(n4), .Z(sum4[3]) );
  CMX2X1 U4 ( .A0(c_out410), .A1(c_out411), .S(n4), .Z(c_out4) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMXI2X1 U7 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CIVX2 U9 ( .A(s43[0]), .Z(n3) );
  CIVX2 U10 ( .A(s44[0]), .Z(n2) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(sum4[2]) );
  CIVX2 U12 ( .A(s43[1]), .Z(n6) );
  CIVX2 U13 ( .A(s44[1]), .Z(n5) );
endmodule


module Add_half_4929 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4930 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2465 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4930 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4929 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4931 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4932 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2466 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4932 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4931 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4933 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4934 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(n1), .B(a), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2467 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_4934 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4933 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4935 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4936 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(n1), .B(a), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2468 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4936 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4935 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_617 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2468 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2467 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2466 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2465 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U4 ( .A(s1), .Z(n3) );
  CIVX1 U5 ( .A(s2), .Z(n2) );
  CMXI2XL U6 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
endmodule


module Add_half_4937 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_4938 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2469 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4938 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4937 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4939 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4940 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2470 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4940 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4939 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4941 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_4942 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX1 U1 ( .A(a), .B(n1), .Z(sum) );
  CIVX2 U2 ( .A(b), .Z(n1) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2471 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_4942 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4941 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4943 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4944 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX1 U1 ( .A(a), .B(n1), .Z(sum) );
  CIVX2 U2 ( .A(b), .Z(n1) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2472 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4944 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4943 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_618 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1;

  Add_full_2472 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2471 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2470 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2469 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_4945 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4946 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2473 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4946 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4945 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4947 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4948 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2474 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4948 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4947 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4949 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4950 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2475 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4950 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4949 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4951 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4952 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2476 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4952 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4951 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_619 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2476 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2475 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2474 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2473 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4953 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4954 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2477 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4954 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4953 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4955 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_4956 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2478 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4956 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4955 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4957 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4958 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2479 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4958 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4957 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4959 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4960 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2480 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4960 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4959 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_620 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2480 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2479 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2478 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2477 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_155 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_620 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_619 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_618 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_617 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n5), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n5), .Z(sum4[0]) );
  CIVX2 U3 ( .A(c_out410), .Z(n3) );
  CMXI2X1 U4 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out4) );
  CIVX2 U5 ( .A(c_out411), .Z(n2) );
  CMX2X1 U6 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2X1 U7 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMXI2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U11 ( .A(n1), .Z(n4) );
  CIVX2 U12 ( .A(c_in4), .Z(n5) );
endmodule


module Add_half_4961 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4962 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2481 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4962 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4961 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4963 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4964 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2482 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4964 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4963 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4965 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4966 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2483 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_4966 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4965 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_4967 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4968 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(n1), .B(a), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2484 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4968 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4967 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_621 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_2484 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2483 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2482 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2481 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CIVX1 U5 ( .A(n2), .Z(n3) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n3), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(c_out10), .A1(c_out11), .S(n3), .Z(c_out2) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_4969 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4970 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2485 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4970 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4969 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4971 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_4972 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2486 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4972 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4971 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_4973 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4974 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2487 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4974 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4973 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_4975 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_4976 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENXL U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2488 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_4976 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4975 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_622 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2488 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2487 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2486 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2485 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2X1 U3 ( .A(c_out00), .B(n1), .Z(n2) );
  CND2X2 U4 ( .A(c_out01), .B(c_in2), .Z(n3) );
  CND2X2 U5 ( .A(n2), .B(n3), .Z(n4) );
  CIVX2 U6 ( .A(c_in2), .Z(n1) );
  CMX2X1 U7 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMX2X1 U9 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_4977 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4978 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2489 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4978 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4977 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4979 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4980 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2490 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4980 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4979 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4981 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4982 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2491 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4982 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4981 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4983 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4984 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2492 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4984 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4983 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_623 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2492 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2491 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2490 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2489 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_4985 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4986 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2493 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4986 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4985 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4987 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4988 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2494 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4988 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4987 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4989 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4990 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2495 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4990 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4989 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4991 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4992 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2496 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4992 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4991 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_624 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2496 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2495 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2494 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2493 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_156 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_624 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_623 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_622 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_621 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n8), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n8), .Z(sum4[0]) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U4 ( .A(c_out411), .Z(n2) );
  CIVX2 U5 ( .A(c_out410), .Z(n3) );
  CIVX1 U6 ( .A(s44[0]), .Z(n4) );
  CIVX1 U7 ( .A(s43[0]), .Z(n5) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(n1), .Z(sum4[2]) );
  CIVX2 U12 ( .A(s43[1]), .Z(n7) );
  CIVX2 U13 ( .A(s44[1]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n1), .Z(sum4[3]) );
  CIVX2 U15 ( .A(c_in4), .Z(n8) );
endmodule


module bit8_39 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n2, n3, n4, n5, n6;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_156 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_155 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_154 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_153 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n6), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n6), .Z(sum8[0]) );
  CMX2X1 U3 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n2) );
  CMX2X2 U4 ( .A0(s83[0]), .A1(s84[0]), .S(n3), .Z(sum8[4]) );
  CIVX1 U5 ( .A(s82[3]), .Z(n4) );
  CMXI2X2 U6 ( .A0(n5), .A1(n4), .S(c_in8), .Z(sum8[3]) );
  CMX2X2 U7 ( .A0(s83[1]), .A1(s84[1]), .S(n2), .Z(sum8[5]) );
  CMX2X2 U8 ( .A0(s83[2]), .A1(s84[2]), .S(n2), .Z(sum8[6]) );
  CMX2X1 U9 ( .A0(s83[3]), .A1(s84[3]), .S(n2), .Z(sum8[7]) );
  CMX2X1 U10 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n3) );
  CMX2X2 U11 ( .A0(c_out810), .A1(c_out811), .S(n3), .Z(c_out8) );
  CMX2X2 U14 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CIVX2 U15 ( .A(s81[3]), .Z(n5) );
  CIVX2 U16 ( .A(c_in8), .Z(n6) );
endmodule


module Add_half_4993 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4994 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2497 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4994 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4993 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4995 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4996 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2498 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4996 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4995 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4997 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_4998 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2499 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_4998 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4997 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_4999 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5000 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2500 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5000 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_4999 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_625 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2500 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2499 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2498 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2497 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5001 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5002 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2501 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5002 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5001 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5003 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5004 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2502 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5004 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5003 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5005 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5006 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2503 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5006 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5005 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5007 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5008 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2504 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5008 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5007 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_626 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2504 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2503 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2502 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2501 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5009 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5010 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2505 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5010 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5009 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5011 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5012 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2506 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5012 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5011 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5013 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5014 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2507 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5014 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5013 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5015 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5016 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2508 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5016 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5015 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_627 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2508 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2507 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2506 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2505 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5017 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5018 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2509 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5018 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5017 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5019 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5020 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2510 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5020 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5019 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5021 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5022 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2511 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5022 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5021 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5023 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5024 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2512 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5024 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5023 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_628 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2512 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2511 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2510 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2509 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_157 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_628 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_627 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_626 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_625 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_5025 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5026 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2513 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5026 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5025 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5027 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5028 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2514 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5028 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5027 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5029 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5030 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2515 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5030 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5029 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5031 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5032 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2516 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5032 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5031 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_629 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2516 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2515 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2514 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2513 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5033 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5034 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2517 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5034 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5033 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5035 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5036 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2518 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5036 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5035 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5037 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5038 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2519 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5038 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5037 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5039 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5040 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2520 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5040 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5039 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_630 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2520 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2519 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2518 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2517 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5041 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5042 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2521 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5042 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5041 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5043 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5044 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2522 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5044 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5043 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5045 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5046 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2523 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5046 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5045 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5047 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5048 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2524 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5048 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5047 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_631 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2524 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2523 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2522 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2521 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5049 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5050 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2525 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5050 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5049 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5051 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5052 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2526 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5052 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5051 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5053 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5054 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2527 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5054 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5053 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5055 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5056 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2528 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5056 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5055 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_632 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2528 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2527 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2526 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2525 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_158 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_632 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_631 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_630 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_629 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_5057 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5058 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2529 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5058 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5057 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5059 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5060 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2530 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5060 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5059 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5061 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5062 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2531 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5062 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5061 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5063 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5064 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2532 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5064 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5063 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_633 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2532 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2531 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2530 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2529 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5065 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5066 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2533 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5066 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5065 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5067 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5068 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2534 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5068 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5067 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5069 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5070 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2535 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5070 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5069 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5071 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5072 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2536 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5072 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5071 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_634 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2536 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2535 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2534 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2533 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5073 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5074 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2537 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5074 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5073 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5075 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5076 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2538 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5076 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5075 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5077 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5078 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2539 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5078 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5077 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5079 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5080 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2540 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5080 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5079 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_635 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2540 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2539 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2538 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2537 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5081 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5082 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2541 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5082 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5081 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5083 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5084 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2542 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5084 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5083 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5085 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5086 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2543 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5086 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5085 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5087 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5088 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2544 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5088 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5087 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_636 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2544 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2543 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2542 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2541 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_159 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_636 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_635 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_634 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_633 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_5089 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5090 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2545 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5090 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5089 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5091 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5092 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2546 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5092 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5091 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5093 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5094 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2547 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5094 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5093 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5095 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5096 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2548 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5096 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5095 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_637 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2548 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2547 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2546 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2545 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5097 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5098 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2549 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5098 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5097 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5099 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5100 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2550 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5100 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5099 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5101 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5102 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2551 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5102 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5101 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5103 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5104 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2552 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5104 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5103 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_638 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2552 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2551 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2550 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2549 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5105 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5106 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2553 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5106 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5105 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5107 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5108 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2554 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5108 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5107 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5109 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5110 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2555 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5110 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5109 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5111 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5112 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2556 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5112 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5111 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_639 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2556 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2555 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2554 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2553 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5113 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5114 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2557 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5114 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5113 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5115 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5116 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2558 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5116 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5115 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5117 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5118 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2559 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5118 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5117 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5119 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5120 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2560 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5120 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5119 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_640 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2560 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2559 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2558 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2557 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_160 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_640 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_639 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_638 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_637 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_40 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n4, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_160 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_159 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_158 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_157 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in8), .Z(n4) );
  CAOR2X1 U6 ( .A(s84[3]), .B(n5), .C(s83[3]), .D(n1), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n5), .C(s83[2]), .D(n1), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n5), .C(s83[1]), .D(n1), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n5), .C(s83[0]), .D(n1), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n4), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n4), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n4), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n4), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n5), .C(c_out810), .D(n1), .Z(c_out8) );
  CANR2X1 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n4), .Z(n1) );
endmodule


module bit32_10 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   c1, c2, c3;

  bit8_40 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8(a32[7:0]), .b8(b32[7:0]), 
        .c_in8(c_in32) );
  bit8_39 A322 ( .sum8(sum32[15:8]), .c_out8(c2), .a8(a32[15:8]), .b8(
        b32[15:8]), .c_in8(c1) );
  bit8_38 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8(a32[23:16]), .b8(
        b32[23:16]), .c_in8(c2) );
  bit8_37 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8(a32[31:24]), .b8(
        b32[31:24]), .c_in8(c3) );
endmodule


module Add_half_5121 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5122 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2561 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5122 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5121 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5123 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5124 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2562 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5124 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5123 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5125 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5126 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2563 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5126 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5125 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5127 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5128 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2564 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5128 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5127 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_641 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2564 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2563 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2562 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2561 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5129 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5130 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2565 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5130 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5129 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5131 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5132 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2566 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5132 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5131 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5133 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5134 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2567 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5134 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5133 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5135 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5136 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2568 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5136 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5135 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_642 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2568 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2567 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2566 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2565 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5137 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5138 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2569 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5138 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5137 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5139 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5140 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2570 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5140 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5139 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5141 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5142 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2571 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5142 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5141 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5143 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5144 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2572 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5144 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5143 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_643 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2572 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2571 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2570 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2569 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5145 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5146 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2573 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5146 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5145 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5147 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5148 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2574 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5148 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5147 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5149 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5150 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2575 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5150 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5149 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5151 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5152 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2576 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5152 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5151 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_644 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2576 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2575 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2574 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2573 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_161 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_644 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_643 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_642 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_641 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_5153 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5154 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2577 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5154 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5153 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5155 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5156 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2578 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5156 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5155 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5157 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5158 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2579 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5158 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5157 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5159 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5160 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2580 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5160 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5159 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_645 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2580 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2579 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2578 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2577 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5161 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5162 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2581 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5162 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5161 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5163 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5164 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2582 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5164 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5163 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5165 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5166 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2583 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5166 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5165 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5167 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5168 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2584 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5168 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5167 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_646 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2584 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2583 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2582 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2581 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5169 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5170 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2585 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5170 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5169 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5171 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5172 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2586 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5172 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5171 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5173 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5174 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2587 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5174 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5173 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5175 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5176 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2588 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5176 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5175 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_647 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2588 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2587 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2586 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2585 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5177 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5178 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2589 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5178 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5177 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5179 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5180 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2590 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5180 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5179 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5181 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5182 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2591 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5182 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5181 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5183 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5184 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2592 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5184 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5183 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_648 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2592 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2591 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2590 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2589 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_162 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_648 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_647 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_646 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_645 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_5185 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5186 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2593 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5186 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5185 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5187 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5188 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2594 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5188 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5187 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5189 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5190 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2595 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5190 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5189 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5191 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5192 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2596 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5192 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5191 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_649 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2596 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2595 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2594 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2593 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5193 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5194 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2597 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5194 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5193 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5195 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5196 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2598 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5196 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5195 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5197 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5198 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2599 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5198 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5197 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5199 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5200 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2600 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5200 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5199 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_650 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2600 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2599 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2598 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2597 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5201 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5202 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2601 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5202 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5201 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5203 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5204 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2602 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5204 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5203 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5205 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5206 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2603 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5206 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5205 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5207 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5208 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2604 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5208 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5207 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_651 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2604 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2603 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2602 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2601 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X2 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CAOR2XL U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
endmodule


module Add_half_5209 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5210 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2605 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5210 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5209 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5211 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5212 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2606 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5212 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5211 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5213 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5214 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2607 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5214 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5213 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5215 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5216 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2608 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5216 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5215 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_652 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2608 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2607 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2606 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2605 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X2 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
endmodule


module bit4_163 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_652 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_651 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_650 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_649 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
endmodule


module Add_half_5217 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5218 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2609 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5218 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5217 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5219 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5220 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2610 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5220 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5219 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5221 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5222 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2611 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5222 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5221 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5223 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5224 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2612 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5224 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5223 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_653 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2612 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2611 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2610 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2609 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5225 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5226 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2613 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5226 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5225 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5227 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5228 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2614 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5228 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5227 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5229 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5230 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2615 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5230 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5229 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5231 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5232 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2616 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5232 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5231 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_654 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2616 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2615 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2614 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2613 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5233 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5234 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2617 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5234 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5233 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5235 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5236 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2618 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5236 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5235 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5237 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5238 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2619 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5238 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5237 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5239 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5240 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2620 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5240 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5239 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_655 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2620 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2619 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2618 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2617 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5241 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5242 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2621 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5242 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5241 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5243 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5244 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2622 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5244 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5243 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5245 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5246 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2623 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5246 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5245 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5247 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5248 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2624 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5248 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5247 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_656 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2624 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2623 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2622 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2621 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_164 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_656 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_655 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_654 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_653 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X2 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2XL U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
endmodule


module bit8_41 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_164 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_163 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_162 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_161 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X2 U3 ( .A0(s83[0]), .A1(s84[0]), .S(n1), .Z(sum8[4]) );
  CMX2X2 U4 ( .A0(s83[1]), .A1(s84[1]), .S(n1), .Z(sum8[5]) );
  CMX2X2 U5 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2X2 U6 ( .A0(s81[0]), .A1(s82[0]), .S(c_in8), .Z(sum8[0]) );
  CMX2X2 U7 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMXI2XL U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out8) );
  CMX2X2 U9 ( .A0(s83[2]), .A1(s84[2]), .S(n1), .Z(sum8[6]) );
  CMX2X2 U10 ( .A0(s83[3]), .A1(s84[3]), .S(n1), .Z(sum8[7]) );
  CMX2X1 U11 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CMX2X1 U12 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CIVX2 U13 ( .A(c_out810), .Z(n3) );
  CIVX2 U14 ( .A(c_out811), .Z(n2) );
endmodule


module Add_half_5249 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5250 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2625 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5250 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5249 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5251 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5252 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2626 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5252 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5251 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5253 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5254 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2627 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5254 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5253 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5255 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5256 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2628 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5256 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5255 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_657 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2628 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2627 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2626 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2625 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_5257 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5258 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2629 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5258 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5257 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5259 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5260 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2630 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5260 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5259 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5261 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5262 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2631 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5262 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5261 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5263 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5264 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2632 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5264 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5263 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_658 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2632 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2631 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2630 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2629 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CIVXL U3 ( .A(s3), .Z(n4) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_5265 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5266 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2633 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5266 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5265 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5267 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5268 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2634 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5268 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5267 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5269 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5270 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2635 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5270 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5269 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5271 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5272 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2636 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5272 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5271 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_659 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2636 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2635 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2634 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2633 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_5273 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5274 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2637 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5274 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5273 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5275 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5276 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2638 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5276 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5275 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5277 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5278 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2639 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5278 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5277 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5279 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5280 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2640 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5280 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5279 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_660 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2640 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2639 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2638 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2637 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX1 U3 ( .A(s3), .Z(n6) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module bit4_165 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_660 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_659 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_658 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_657 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n5), .Z(sum4[0]) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
  CIVX2 U12 ( .A(c_in4), .Z(n5) );
endmodule


module Add_half_5281 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5282 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2641 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5282 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5281 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5283 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5284 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2642 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5284 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5283 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5285 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5286 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2643 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5286 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5285 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5287 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5288 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2644 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5288 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5287 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_661 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2644 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2643 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2642 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2641 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_5289 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5290 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2645 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5290 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5289 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5291 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5292 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2646 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5292 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5291 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5293 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5294 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2647 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5294 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5293 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5295 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5296 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2648 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5296 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5295 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_662 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2648 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2647 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2646 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2645 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5297 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5298 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2649 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5298 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5297 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5299 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5300 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2650 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5300 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5299 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5301 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5302 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2651 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5302 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5301 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5303 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5304 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2652 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5304 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5303 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_663 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2652 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2651 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2650 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2649 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_5305 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5306 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2653 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5306 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5305 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5307 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5308 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2654 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5308 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5307 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5309 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5310 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2655 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5310 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5309 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5311 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5312 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2656 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5312 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5311 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_664 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2656 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2655 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2654 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2653 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module bit4_166 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_664 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_663 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_662 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_661 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n11), .Z(sum4[0]) );
  CIVX2 U3 ( .A(c_out410), .Z(n3) );
  CIVX2 U4 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n8) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U8 ( .A(s41[1]), .Z(n5) );
  CIVX2 U10 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(s43[0]), .Z(n7) );
  CIVX2 U13 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX2 U15 ( .A(s43[1]), .Z(n10) );
  CIVX2 U16 ( .A(s44[1]), .Z(n9) );
  CMXI2X1 U17 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
  CIVX2 U18 ( .A(c_in4), .Z(n11) );
endmodule


module Add_half_5313 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5314 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2657 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5314 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5313 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5315 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5316 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2658 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5316 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5315 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5317 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5318 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2659 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5318 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5317 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5319 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5320 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2660 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5320 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5319 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_665 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2660 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2659 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2658 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2657 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(n1), .Z(n2) );
  CIVX2 U6 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_5321 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5322 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2661 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5322 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5321 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5323 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5324 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2662 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5324 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5323 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5325 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5326 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2663 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5326 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5325 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5327 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5328 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2664 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5328 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5327 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_666 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2664 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2663 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2662 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2661 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVXL U5 ( .A(s3), .Z(n3) );
  CMX2X1 U6 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CIVX2 U8 ( .A(s4), .Z(n2) );
  CIVX2 U9 ( .A(c_in2), .Z(n4) );
endmodule


module Add_half_5329 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5330 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2665 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5330 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5329 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5331 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5332 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2666 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5332 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5331 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5333 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5334 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2667 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5334 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5333 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5335 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5336 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2668 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5336 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5335 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_667 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_2668 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2667 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2666 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2665 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_5337 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5338 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2669 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5338 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5337 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5339 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5340 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2670 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5340 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5339 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5341 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_5342 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2671 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5342 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5341 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5343 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5344 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2672 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5344 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5343 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_668 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2672 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2671 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2670 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2669 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(s3), .Z(n6) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module bit4_167 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_668 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_667 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_666 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_665 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module Add_half_5345 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5346 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2673 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5346 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5345 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5347 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5348 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2674 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5348 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5347 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5349 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5350 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2675 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5350 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5349 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5351 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5352 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2676 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5352 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5351 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_669 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_2676 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2675 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2674 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2673 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n3), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(c_in2), .Z(n3) );
endmodule


module Add_half_5353 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5354 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2677 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5354 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5353 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5355 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5356 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2678 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5356 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5355 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5357 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5358 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2679 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5358 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5357 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5359 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5360 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2680 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5360 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5359 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_670 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_2680 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2679 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2678 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2677 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n2), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CIVX2 U6 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_5361 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5362 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2681 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5362 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5361 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5363 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5364 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2682 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5364 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5363 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5365 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5366 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2683 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5366 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5365 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5367 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5368 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2684 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5368 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5367 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_671 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2684 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2683 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2682 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2681 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_5369 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5370 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2685 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5370 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5369 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5371 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5372 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2686 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5372 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5371 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5373 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5374 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2687 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5374 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5373 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5375 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5376 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2688 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5376 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5375 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_672 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2688 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2687 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2686 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2685 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_168 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_672 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_671 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_670 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_669 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(c_out410), .Z(n3) );
  CIVX2 U4 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n10) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n10), .Z(c_out4) );
  CIVX2 U8 ( .A(s41[0]), .Z(n5) );
  CIVX2 U9 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U11 ( .A(s41[1]), .Z(n7) );
  CIVX2 U12 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U13 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n9) );
  CIVX2 U15 ( .A(s44[0]), .Z(n8) );
  CMXI2X1 U16 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CIVX2 U17 ( .A(s43[1]), .Z(n12) );
  CIVX2 U18 ( .A(s44[1]), .Z(n11) );
  CMXI2X1 U19 ( .A0(n12), .A1(n11), .S(n10), .Z(sum4[3]) );
endmodule


module bit8_42 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_168 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_167 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_166 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_165 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X2 U3 ( .A0(s83[2]), .A1(s84[2]), .S(n9), .Z(sum8[6]) );
  CMX2X2 U4 ( .A0(s83[1]), .A1(s84[1]), .S(n1), .Z(sum8[5]) );
  CIVXL U5 ( .A(n10), .Z(n1) );
  CND2X1 U6 ( .A(s83[0]), .B(n2), .Z(n3) );
  CND2X1 U7 ( .A(s84[0]), .B(n8), .Z(n4) );
  CND2X4 U8 ( .A(n3), .B(n4), .Z(sum8[4]) );
  CIVXL U9 ( .A(n8), .Z(n2) );
  CIVX2 U10 ( .A(n10), .Z(n8) );
  CND2X1 U11 ( .A(s81[0]), .B(n5), .Z(n6) );
  CND2X1 U12 ( .A(s82[0]), .B(c_in8), .Z(n7) );
  CND2X4 U13 ( .A(n6), .B(n7), .Z(sum8[0]) );
  CIVXL U14 ( .A(c_in8), .Z(n5) );
  CMX2X2 U15 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMXI2X1 U16 ( .A0(n12), .A1(n11), .S(n8), .Z(c_out8) );
  CMX2XL U17 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n9) );
  CMX2X1 U18 ( .A0(s83[3]), .A1(s84[3]), .S(n9), .Z(sum8[7]) );
  CMX2X1 U19 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2X1 U20 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CIVX2 U21 ( .A(c_out810), .Z(n12) );
  CIVX2 U22 ( .A(c_out811), .Z(n11) );
  CMXI2X1 U23 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n10) );
endmodule


module Add_half_5377 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5378 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2689 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5378 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5377 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5379 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5380 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2690 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5380 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5379 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5381 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5382 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2691 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5382 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5381 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5383 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5384 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2692 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5384 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5383 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_673 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2692 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2691 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2690 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2689 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVXL U3 ( .A(s3), .Z(n6) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CIVX2 U7 ( .A(s1), .Z(n3) );
  CIVX2 U8 ( .A(s2), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_5385 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5386 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2693 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5386 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5385 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5387 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5388 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2694 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5388 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5387 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5389 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_5390 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2695 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5390 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5389 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5391 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5392 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2696 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5392 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5391 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_674 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2696 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2695 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2694 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2693 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U7 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_5393 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5394 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2697 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5394 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5393 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5395 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5396 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2698 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5396 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5395 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5397 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5398 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2699 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5398 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5397 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5399 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5400 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2700 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5400 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5399 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_675 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_2700 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2699 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2698 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2697 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_5401 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_5402 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2701 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5402 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5401 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5403 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5404 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2702 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5404 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5403 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5405 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_5406 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2703 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5406 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5405 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5407 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5408 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2704 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5408 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5407 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_676 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2704 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2703 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2702 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2701 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_169 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_676 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_675 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_674 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_673 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2XL U4 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module Add_half_5409 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5410 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2705 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5410 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5409 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5411 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5412 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2706 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5412 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5411 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5413 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5414 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2707 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5414 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5413 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5415 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5416 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2708 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5416 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5415 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_677 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2708 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2707 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2706 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2705 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_5417 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5418 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2709 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5418 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5417 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5419 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5420 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2710 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5420 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5419 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5421 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5422 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2711 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5422 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5421 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5423 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5424 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2712 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5424 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5423 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_678 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_2712 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2711 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2710 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2709 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_5425 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5426 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2713 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5426 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5425 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5427 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5428 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2714 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5428 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5427 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5429 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5430 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2715 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5430 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5429 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5431 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5432 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2716 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5432 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5431 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_679 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2716 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2715 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2714 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2713 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U4 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMX2XL U5 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n4) );
  CIVX2 U8 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
endmodule


module Add_half_5433 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5434 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2717 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5434 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5433 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5435 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5436 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2718 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5436 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5435 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5437 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5438 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2719 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5438 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5437 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5439 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5440 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2720 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5440 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5439 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_680 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2720 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2719 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2718 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2717 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_170 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_680 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_679 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_678 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_677 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(c_out410), .A1(c_out411), .S(n8), .Z(c_out4) );
  CMXI2X1 U4 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U5 ( .A(n1), .Z(n8) );
  CIVX2 U6 ( .A(s41[0]), .Z(n3) );
  CIVX2 U7 ( .A(s42[0]), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U9 ( .A(s41[1]), .Z(n5) );
  CIVX2 U10 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(s43[0]), .Z(n7) );
  CIVX2 U13 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX2 U15 ( .A(s43[1]), .Z(n10) );
  CIVX2 U16 ( .A(s44[1]), .Z(n9) );
  CMXI2X1 U17 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
endmodule


module Add_half_5441 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5442 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2721 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5442 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5441 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5443 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5444 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2722 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5444 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5443 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5445 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5446 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2723 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5446 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5445 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5447 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5448 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2724 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5448 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5447 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_681 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2724 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2723 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2722 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2721 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CIVX2 U4 ( .A(c_in2), .Z(n2) );
  CMXI2XL U5 ( .A0(n6), .A1(n5), .S(n1), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CIVX2 U7 ( .A(s1), .Z(n4) );
  CIVX2 U8 ( .A(s2), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module Add_half_5449 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_5450 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2725 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5450 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5449 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5451 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5452 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2726 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5452 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5451 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5453 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_5454 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2727 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5454 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5453 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5455 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5456 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2728 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5456 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5455 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_682 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_2728 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2727 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2726 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2725 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_5457 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_5458 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2729 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5458 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5457 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5459 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5460 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2730 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5460 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5459 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5461 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5462 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2731 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5462 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5461 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_5463 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5464 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2732 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5464 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5463 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_683 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2732 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2731 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2730 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2729 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U4 ( .A(s2), .Z(n5) );
  CIVX1 U5 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U6 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CIVXL U7 ( .A(s1), .Z(n6) );
  CMX2XL U8 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CIVX2 U9 ( .A(c_out10), .Z(n4) );
  CMXI2X1 U10 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_5465 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5466 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2733 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5466 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5465 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5467 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5468 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2734 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5468 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5467 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5469 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_5470 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2735 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5470 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5469 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5471 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5472 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX1 U1 ( .A(a), .B(n1), .Z(sum) );
  CIVX20 U2 ( .A(b), .Z(n1) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2736 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5472 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5471 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_684 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2736 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2735 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2734 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2733 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n2) );
  CIVX1 U4 ( .A(c_out10), .Z(n5) );
  CMX2XL U5 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CIVX1 U6 ( .A(c_out11), .Z(n4) );
  CMXI2X1 U7 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CMXI2X1 U8 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n3) );
  CMXI2XL U9 ( .A0(n7), .A1(n6), .S(n1), .Z(sum2[1]) );
  CMX2X1 U10 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n7) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
endmodule


module bit4_171 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_684 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_683 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_682 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_681 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMX2XL U4 ( .A0(s44[0]), .A1(s43[0]), .S(n1), .Z(sum4[2]) );
  CIVX1 U5 ( .A(c_out411), .Z(n2) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMX2XL U7 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2X1 U8 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U9 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U10 ( .A(c_out410), .Z(n3) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module Add_half_5473 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5474 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2737 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5474 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5473 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5475 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5476 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2738 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5476 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5475 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5477 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5478 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2739 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5478 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5477 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5479 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5480 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2740 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5480 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5479 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_685 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_2740 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2739 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2738 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2737 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_5481 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5482 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2741 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5482 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5481 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5483 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5484 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2742 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5484 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5483 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5485 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5486 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2743 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5486 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5485 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5487 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5488 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2744 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5488 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5487 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_686 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_2744 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2743 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2742 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2741 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_5489 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_5490 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2745 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5490 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5489 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5491 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5492 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2746 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5492 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5491 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5493 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5494 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2747 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5494 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5493 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5495 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5496 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2748 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5496 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5495 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_687 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2748 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2747 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2746 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2745 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_5497 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_5498 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2749 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5498 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5497 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5499 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5500 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2750 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5500 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5499 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5501 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5502 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2751 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5502 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5501 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5503 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X2 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5504 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2752 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5504 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5503 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_688 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2752 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2751 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2750 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2749 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_172 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_688 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_687 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_686 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_685 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVXL U3 ( .A(n10), .Z(n1) );
  CIVXL U4 ( .A(n1), .Z(n2) );
  CIVX1 U5 ( .A(s41[0]), .Z(n7) );
  CIVX1 U6 ( .A(c_out410), .Z(n5) );
  CMXI2XL U7 ( .A0(n12), .A1(n11), .S(n2), .Z(sum4[3]) );
  CMX2X1 U8 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U9 ( .A(c_out411), .Z(n4) );
  CMXI2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n3) );
  CIVX2 U11 ( .A(n3), .Z(n10) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(n10), .Z(c_out4) );
  CIVX2 U13 ( .A(s42[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U15 ( .A(s43[0]), .Z(n9) );
  CIVX2 U16 ( .A(s44[0]), .Z(n8) );
  CMXI2X1 U17 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CIVX2 U18 ( .A(s43[1]), .Z(n12) );
  CIVX2 U19 ( .A(s44[1]), .Z(n11) );
endmodule


module bit8_43 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_172 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_171 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_170 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_169 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVX3 U3 ( .A(n2), .Z(sum8[4]) );
  CIVX2 U4 ( .A(n1), .Z(c_out8) );
  CMXI2X2 U5 ( .A0(n10), .A1(n9), .S(c_in8), .Z(sum8[0]) );
  CMXI2X1 U6 ( .A0(c_out810), .A1(c_out811), .S(n8), .Z(n1) );
  CMXI2X1 U7 ( .A0(s83[0]), .A1(s84[0]), .S(n8), .Z(n2) );
  CIVX1 U8 ( .A(s84[3]), .Z(n15) );
  CIVX1 U9 ( .A(n8), .Z(n3) );
  CIVX2 U10 ( .A(n3), .Z(n4) );
  CIVXL U11 ( .A(s82[2]), .Z(n13) );
  CMX2X1 U12 ( .A0(s83[1]), .A1(s84[1]), .S(n8), .Z(sum8[5]) );
  CND2X1 U13 ( .A(c_out800), .B(n5), .Z(n6) );
  CND2X1 U14 ( .A(c_out801), .B(c_in8), .Z(n7) );
  CND2X2 U15 ( .A(n6), .B(n7), .Z(n8) );
  CIVX2 U16 ( .A(c_in8), .Z(n5) );
  CMXI2X1 U17 ( .A0(n14), .A1(n13), .S(c_in8), .Z(sum8[2]) );
  CMX2X2 U18 ( .A0(s83[2]), .A1(s84[2]), .S(n4), .Z(sum8[6]) );
  CMX2X2 U19 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CIVX1 U20 ( .A(s82[1]), .Z(n11) );
  CIVX1 U21 ( .A(s82[0]), .Z(n9) );
  CIVX1 U22 ( .A(s81[0]), .Z(n10) );
  CMXI2X2 U23 ( .A0(n16), .A1(n15), .S(n4), .Z(sum8[7]) );
  CIVX1 U24 ( .A(s81[2]), .Z(n14) );
  CIVX2 U25 ( .A(s81[1]), .Z(n12) );
  CMXI2X1 U26 ( .A0(n12), .A1(n11), .S(c_in8), .Z(sum8[1]) );
  CIVX2 U27 ( .A(s83[3]), .Z(n16) );
endmodule


module Add_half_5505 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5506 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2753 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5506 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5505 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5507 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5508 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2754 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5508 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5507 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5509 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5510 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2755 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5510 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5509 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5511 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5512 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2756 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5512 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5511 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_689 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2756 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2755 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2754 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2753 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5513 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5514 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2757 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5514 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5513 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5515 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5516 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2758 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5516 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5515 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5517 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5518 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2759 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5518 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5517 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5519 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5520 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2760 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5520 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5519 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_690 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2760 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2759 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2758 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2757 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5521 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5522 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2761 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5522 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5521 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5523 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5524 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2762 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5524 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5523 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5525 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5526 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2763 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5526 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5525 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5527 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5528 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2764 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5528 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5527 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_691 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2764 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2763 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2762 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2761 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5529 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5530 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2765 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5530 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5529 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5531 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5532 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2766 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5532 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5531 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5533 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5534 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2767 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5534 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5533 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5535 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5536 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2768 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5536 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5535 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_692 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2768 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2767 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2766 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2765 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_173 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_692 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_691 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_690 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_689 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_5537 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5538 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2769 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5538 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5537 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5539 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5540 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2770 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5540 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5539 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5541 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5542 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2771 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5542 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5541 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5543 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5544 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2772 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5544 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5543 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_693 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2772 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2771 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2770 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2769 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5545 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5546 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2773 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5546 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5545 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5547 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5548 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2774 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5548 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5547 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5549 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5550 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2775 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5550 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5549 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5551 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5552 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2776 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5552 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5551 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_694 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2776 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2775 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2774 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2773 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5553 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5554 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2777 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5554 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5553 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5555 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5556 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2778 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5556 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5555 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5557 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5558 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2779 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5558 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5557 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5559 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5560 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2780 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5560 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5559 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_695 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2780 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2779 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2778 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2777 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5561 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5562 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2781 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5562 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5561 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5563 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5564 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2782 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5564 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5563 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5565 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5566 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2783 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5566 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5565 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5567 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5568 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2784 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5568 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5567 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_696 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2784 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2783 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2782 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2781 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_174 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_696 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_695 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_694 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_693 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_5569 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5570 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2785 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5570 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5569 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5571 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5572 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2786 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5572 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5571 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5573 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5574 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2787 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5574 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5573 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5575 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5576 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2788 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5576 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5575 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_697 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2788 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2787 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2786 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2785 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5577 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5578 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2789 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5578 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5577 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5579 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5580 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2790 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5580 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5579 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5581 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5582 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2791 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5582 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5581 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5583 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5584 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2792 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5584 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5583 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_698 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2792 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2791 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2790 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2789 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5585 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5586 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2793 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5586 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5585 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5587 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5588 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2794 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5588 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5587 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5589 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5590 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2795 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5590 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5589 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5591 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5592 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2796 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5592 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5591 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_699 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2796 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2795 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2794 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2793 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5593 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5594 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2797 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5594 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5593 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5595 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5596 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2798 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5596 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5595 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5597 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5598 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2799 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5598 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5597 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5599 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5600 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2800 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5600 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5599 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_700 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2800 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2799 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2798 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2797 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_175 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_700 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_699 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_698 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_697 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_5601 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5602 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2801 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5602 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5601 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5603 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5604 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2802 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5604 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5603 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5605 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5606 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2803 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5606 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5605 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5607 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5608 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2804 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5608 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5607 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_701 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2804 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2803 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2802 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2801 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5609 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5610 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2805 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5610 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5609 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5611 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5612 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2806 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5612 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5611 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5613 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5614 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2807 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5614 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5613 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5615 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5616 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2808 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5616 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5615 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_702 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2808 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2807 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2806 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2805 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5617 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5618 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2809 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5618 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5617 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5619 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5620 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2810 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5620 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5619 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5621 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5622 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2811 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5622 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5621 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5623 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5624 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2812 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5624 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5623 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_703 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2812 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2811 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2810 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2809 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5625 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5626 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2813 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5626 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5625 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5627 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5628 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2814 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5628 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5627 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5629 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5630 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2815 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5630 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5629 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5631 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5632 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2816 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5632 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5631 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_704 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2816 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2815 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2814 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2813 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_176 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_704 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_703 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_702 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_701 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_44 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n4, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_176 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_175 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_174 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_173 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in8), .Z(n4) );
  CAOR2X1 U6 ( .A(s84[3]), .B(n5), .C(s83[3]), .D(n1), .Z(sum8[7]) );
  CAOR2X1 U7 ( .A(s84[2]), .B(n5), .C(s83[2]), .D(n1), .Z(sum8[6]) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n5), .C(s83[1]), .D(n1), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n5), .C(s83[0]), .D(n1), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n4), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n4), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n4), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n4), .Z(sum8[0]) );
  CAOR2X1 U14 ( .A(c_out811), .B(n5), .C(c_out810), .D(n1), .Z(c_out8) );
  CANR2X1 U3 ( .A(c_out801), .B(c_in8), .C(c_out800), .D(n4), .Z(n1) );
endmodule


module bit32_11 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   c1, c2, c3, n1, n2;

  bit8_44 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8(a32[7:0]), .b8(b32[7:0]), 
        .c_in8(c_in32) );
  bit8_43 A322 ( .sum8(sum32[15:8]), .c_out8(c2), .a8(a32[15:8]), .b8(
        b32[15:8]), .c_in8(c1) );
  bit8_42 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8(a32[23:16]), .b8(
        b32[23:16]), .c_in8(c2) );
  bit8_41 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8(a32[31:24]), .b8(
        b32[31:24]), .c_in8(n2) );
  CIVX1 U1 ( .A(c3), .Z(n1) );
  CIVX3 U2 ( .A(n1), .Z(n2) );
endmodule


module Add_half_5633 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5634 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2817 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5634 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5633 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5635 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5636 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2818 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5636 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5635 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5637 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5638 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2819 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5638 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5637 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5639 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5640 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2820 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5640 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5639 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_705 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2820 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2819 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2818 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2817 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5641 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5642 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2821 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5642 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5641 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5643 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5644 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2822 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5644 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5643 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5645 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5646 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2823 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5646 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5645 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5647 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5648 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2824 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5648 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5647 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_706 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2824 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2823 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2822 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2821 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5649 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5650 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2825 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5650 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5649 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5651 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5652 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2826 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5652 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5651 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5653 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5654 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2827 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5654 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5653 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5655 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5656 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2828 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5656 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5655 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_707 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2828 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2827 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2826 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2825 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5657 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5658 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2829 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5658 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5657 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5659 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5660 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2830 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5660 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5659 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5661 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5662 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2831 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5662 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5661 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5663 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5664 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2832 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5664 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5663 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_708 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2832 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2831 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2830 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2829 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_177 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_708 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_707 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_706 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_705 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_5665 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5666 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2833 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5666 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5665 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5667 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5668 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2834 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5668 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5667 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5669 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5670 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2835 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5670 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5669 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5671 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5672 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2836 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5672 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5671 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_709 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2836 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2835 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2834 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2833 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5673 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5674 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2837 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5674 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5673 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5675 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5676 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2838 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5676 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5675 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5677 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5678 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2839 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5678 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5677 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5679 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5680 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2840 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5680 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5679 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_710 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2840 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2839 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2838 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2837 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5681 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5682 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2841 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5682 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5681 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5683 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5684 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2842 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5684 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5683 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5685 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5686 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2843 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5686 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5685 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5687 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5688 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2844 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5688 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5687 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_711 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2844 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2843 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2842 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2841 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5689 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5690 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2845 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5690 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5689 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5691 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5692 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2846 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5692 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5691 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5693 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5694 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2847 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5694 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5693 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5695 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5696 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2848 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5696 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5695 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_712 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2848 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2847 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2846 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2845 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_178 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_712 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_711 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_710 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_709 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_5697 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5698 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2849 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5698 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5697 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5699 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5700 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2850 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5700 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5699 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5701 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5702 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2851 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5702 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5701 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5703 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5704 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2852 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5704 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5703 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_713 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2852 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2851 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2850 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2849 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5705 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5706 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2853 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5706 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5705 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5707 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5708 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2854 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5708 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5707 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5709 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5710 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2855 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5710 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5709 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5711 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5712 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2856 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5712 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5711 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_714 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2856 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2855 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2854 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2853 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5713 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5714 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2857 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5714 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5713 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5715 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5716 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2858 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5716 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5715 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5717 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5718 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2859 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5718 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5717 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5719 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5720 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2860 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5720 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5719 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_715 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2860 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2859 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2858 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2857 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5721 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5722 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2861 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5722 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5721 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5723 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5724 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2862 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5724 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5723 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5725 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5726 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2863 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5726 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5725 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5727 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5728 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2864 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5728 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5727 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_716 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2864 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2863 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2862 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2861 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_179 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_716 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_715 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_714 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_713 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_5729 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5730 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2865 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5730 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5729 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5731 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5732 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2866 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5732 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5731 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5733 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5734 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2867 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5734 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5733 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5735 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5736 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2868 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5736 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5735 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_717 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2868 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2867 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2866 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2865 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5737 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5738 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2869 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5738 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5737 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5739 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5740 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2870 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5740 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5739 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5741 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5742 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2871 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5742 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5741 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5743 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5744 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2872 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5744 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5743 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_718 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2872 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2871 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2870 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2869 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5745 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5746 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2873 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5746 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5745 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5747 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5748 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2874 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5748 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5747 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5749 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5750 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2875 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5750 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5749 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5751 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5752 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2876 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5752 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5751 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_719 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2876 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2875 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2874 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2873 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5753 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5754 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2877 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5754 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5753 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5755 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5756 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2878 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5756 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5755 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5757 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5758 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2879 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5758 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5757 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5759 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5760 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2880 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5760 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5759 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_720 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2880 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2879 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2878 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2877 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_180 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_720 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_719 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_718 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_717 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_45 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_180 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_179 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_178 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_177 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out8) );
  CMX2X1 U4 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CMXI2X4 U5 ( .A0(n5), .A1(n4), .S(c_in8), .Z(sum8[0]) );
  CMX2XL U6 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2X1 U7 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2XL U8 ( .A0(s83[3]), .A1(s84[3]), .S(n1), .Z(sum8[7]) );
  CMX2X2 U9 ( .A0(s83[0]), .A1(s84[0]), .S(n1), .Z(sum8[4]) );
  CMX2X1 U10 ( .A0(s83[2]), .A1(s84[2]), .S(n1), .Z(sum8[6]) );
  CMX2X1 U11 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2X1 U12 ( .A0(s83[1]), .A1(s84[1]), .S(n1), .Z(sum8[5]) );
  CIVX2 U13 ( .A(c_out810), .Z(n3) );
  CIVX2 U14 ( .A(c_out811), .Z(n2) );
  CIVX2 U15 ( .A(s81[0]), .Z(n5) );
  CIVX2 U16 ( .A(s82[0]), .Z(n4) );
endmodule


module Add_half_5761 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5762 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2881 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5762 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5761 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5763 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5764 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2882 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5764 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5763 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5765 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5766 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2883 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5766 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5765 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5767 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5768 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2884 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5768 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5767 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_721 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2884 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2883 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2882 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2881 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_5769 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5770 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2885 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5770 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5769 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5771 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5772 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2886 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5772 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5771 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5773 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5774 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2887 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5774 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5773 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5775 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5776 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2888 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5776 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5775 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_722 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2888 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2887 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2886 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2885 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_5777 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5778 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2889 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5778 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5777 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5779 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5780 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2890 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5780 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5779 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5781 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5782 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2891 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5782 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5781 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5783 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5784 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2892 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5784 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5783 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_723 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2892 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2891 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2890 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2889 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_5785 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5786 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2893 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5786 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5785 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5787 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5788 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2894 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5788 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5787 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5789 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5790 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2895 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5790 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5789 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5791 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5792 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2896 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5792 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5791 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_724 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2896 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2895 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2894 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2893 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVXL U3 ( .A(s3), .Z(n6) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module bit4_181 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_724 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_723 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_722 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_721 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n5), .Z(sum4[0]) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
  CIVX2 U12 ( .A(c_in4), .Z(n5) );
endmodule


module Add_half_5793 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5794 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2897 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5794 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5793 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5795 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5796 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2898 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5796 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5795 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5797 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5798 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2899 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5798 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5797 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5799 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5800 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2900 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5800 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5799 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_725 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2900 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2899 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2898 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2897 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_5801 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5802 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2901 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5802 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5801 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5803 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_5804 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2902 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5804 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5803 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5805 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5806 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_2903 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5806 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5805 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5807 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5808 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2904 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5808 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5807 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_726 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_2904 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2903 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2902 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2901 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_5809 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5810 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2905 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5810 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5809 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5811 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5812 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2906 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5812 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5811 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_5813 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5814 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2907 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5814 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5813 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_5815 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5816 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2908 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5816 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5815 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_727 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2908 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2907 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2906 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2905 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_5817 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5818 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2909 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5818 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5817 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5819 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5820 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_2910 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5820 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5819 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5821 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5822 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2911 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5822 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5821 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5823 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5824 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2912 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5824 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5823 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_728 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2912 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2911 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2910 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2909 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module bit4_182 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_728 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_727 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_726 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_725 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n11), .Z(sum4[0]) );
  CIVX2 U3 ( .A(c_out410), .Z(n3) );
  CIVX2 U4 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n8) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U8 ( .A(s41[1]), .Z(n5) );
  CIVX2 U10 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(s43[0]), .Z(n7) );
  CIVX2 U13 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX2 U15 ( .A(s43[1]), .Z(n10) );
  CIVX2 U16 ( .A(s44[1]), .Z(n9) );
  CMXI2X1 U17 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
  CIVX2 U18 ( .A(c_in4), .Z(n11) );
endmodule


module Add_half_5825 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5826 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2913 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5826 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5825 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5827 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5828 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2914 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5828 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5827 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5829 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5830 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2915 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5830 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5829 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5831 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5832 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2916 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5832 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5831 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_729 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2916 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2915 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2914 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2913 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_5833 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5834 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2917 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5834 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5833 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5835 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5836 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2918 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5836 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5835 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5837 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5838 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2919 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5838 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5837 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5839 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5840 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2920 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5840 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5839 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_730 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_2920 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2919 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2918 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2917 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_5841 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5842 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2921 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5842 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5841 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5843 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5844 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2922 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5844 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5843 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5845 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5846 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2923 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5846 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5845 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5847 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5848 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2924 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5848 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5847 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_731 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_2924 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2923 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2922 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2921 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_5849 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5850 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2925 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5850 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5849 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5851 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5852 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2926 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5852 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5851 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5853 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_5854 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2927 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5854 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5853 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5855 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5856 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2928 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5856 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5855 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_732 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2928 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2927 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2926 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2925 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s3), .Z(n6) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module bit4_183 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_732 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_731 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_730 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_729 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2X1 U4 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U6 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module Add_half_5857 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5858 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2929 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5858 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5857 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5859 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5860 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2930 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5860 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5859 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5861 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5862 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2931 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5862 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5861 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5863 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5864 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2932 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5864 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5863 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_733 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2932 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2931 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2930 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2929 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_5865 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5866 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2933 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5866 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5865 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5867 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5868 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2934 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5868 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5867 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5869 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5870 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2935 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5870 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5869 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5871 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5872 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2936 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5872 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5871 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_734 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2936 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2935 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2934 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2933 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_5873 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5874 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2937 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5874 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5873 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5875 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5876 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2938 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5876 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5875 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5877 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5878 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2939 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5878 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5877 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5879 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5880 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2940 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5880 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5879 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_735 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2940 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2939 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2938 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2937 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_5881 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5882 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2941 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5882 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5881 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5883 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5884 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2942 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5884 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5883 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5885 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5886 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2943 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5886 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5885 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5887 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5888 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2944 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5888 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5887 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_736 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2944 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2943 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2942 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2941 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_184 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_736 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_735 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_734 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_733 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n10), .Z(c_out4) );
  CIVX2 U4 ( .A(c_out410), .Z(n3) );
  CIVX2 U5 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n10) );
  CIVX2 U8 ( .A(s41[0]), .Z(n5) );
  CIVX2 U9 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U11 ( .A(s41[1]), .Z(n7) );
  CIVX2 U12 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U13 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n9) );
  CIVX2 U15 ( .A(s44[0]), .Z(n8) );
  CMXI2X1 U16 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CIVX2 U17 ( .A(s43[1]), .Z(n12) );
  CIVX2 U18 ( .A(s44[1]), .Z(n11) );
  CMXI2X1 U19 ( .A0(n12), .A1(n11), .S(n10), .Z(sum4[3]) );
endmodule


module bit8_46 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   n14, c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n6, n7,
         n8, n9, n10, n11, n12, n13;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_184 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_183 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_182 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_181 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CIVX2 U3 ( .A(n6), .Z(n13) );
  CMXI2X1 U4 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CMXI2X2 U5 ( .A0(n9), .A1(n10), .S(n3), .Z(sum8[3]) );
  CMX2X1 U6 ( .A0(s83[3]), .A1(s84[3]), .S(n2), .Z(sum8[7]) );
  CMX2X2 U7 ( .A0(s83[1]), .A1(s84[1]), .S(n2), .Z(sum8[5]) );
  CIVX1 U8 ( .A(n1), .Z(n2) );
  CMX2X2 U9 ( .A0(s83[2]), .A1(s84[2]), .S(n2), .Z(sum8[6]) );
  CIVXL U10 ( .A(c_in8), .Z(n3) );
  CIVX2 U11 ( .A(n14), .Z(n4) );
  CIVX4 U12 ( .A(n4), .Z(sum8[4]) );
  CMXI2X1 U13 ( .A0(n12), .A1(n11), .S(n13), .Z(n14) );
  CMX2X2 U14 ( .A0(s81[0]), .A1(s82[0]), .S(c_in8), .Z(sum8[0]) );
  CMX2X2 U15 ( .A0(c_out810), .A1(c_out811), .S(n13), .Z(c_out8) );
  CMX2X1 U16 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMXI2X2 U17 ( .A0(n8), .A1(n7), .S(c_in8), .Z(sum8[2]) );
  CMXI2X1 U18 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n6) );
  CIVX2 U19 ( .A(s81[2]), .Z(n8) );
  CIVX2 U20 ( .A(s82[2]), .Z(n7) );
  CIVX2 U21 ( .A(s81[3]), .Z(n10) );
  CIVX2 U22 ( .A(s82[3]), .Z(n9) );
  CIVX2 U23 ( .A(s83[0]), .Z(n12) );
  CIVX2 U24 ( .A(s84[0]), .Z(n11) );
endmodule


module Add_half_5889 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5890 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2945 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5890 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5889 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5891 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5892 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2946 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5892 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5891 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5893 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5894 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2947 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5894 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5893 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5895 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5896 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2948 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5896 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5895 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_737 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2948 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2947 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2946 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2945 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_5897 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5898 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2949 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5898 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5897 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5899 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5900 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2950 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5900 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5899 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5901 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_5902 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2951 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5902 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5901 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5903 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5904 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2952 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5904 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5903 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_738 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2952 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2951 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2950 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2949 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX1 U4 ( .A(c_out10), .Z(n3) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_5905 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5906 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2953 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5906 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5905 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5907 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5908 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2954 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5908 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5907 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5909 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5910 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2955 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5910 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5909 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5911 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5912 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2956 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5912 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5911 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_739 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2956 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2955 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2954 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2953 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_5913 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5914 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2957 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5914 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5913 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5915 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5916 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2958 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5916 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5915 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5917 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_5918 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2959 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5918 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5917 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5919 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5920 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2960 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5920 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5919 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_740 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2960 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2959 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2958 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2957 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_185 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_740 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_739 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_738 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_737 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U4 ( .A0(c_out410), .A1(c_out411), .S(n4), .Z(c_out4) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CIVX2 U8 ( .A(s41[1]), .Z(n3) );
  CIVX2 U9 ( .A(s42[1]), .Z(n2) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U11 ( .A(s43[1]), .Z(n6) );
  CIVX2 U12 ( .A(s44[1]), .Z(n5) );
  CMXI2X1 U13 ( .A0(n6), .A1(n5), .S(n4), .Z(sum4[3]) );
endmodule


module Add_half_5921 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5922 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2961 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5922 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5921 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5923 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5924 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2962 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5924 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5923 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5925 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5926 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2963 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5926 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5925 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5927 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5928 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2964 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5928 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5927 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_741 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2964 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2963 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2962 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2961 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(n1), .Z(n4) );
  CIVX2 U6 ( .A(s1), .Z(n3) );
  CIVX2 U7 ( .A(s2), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_5929 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5930 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2965 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5930 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5929 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5931 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5932 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2966 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5932 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5931 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5933 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_5934 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2967 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5934 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5933 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5935 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5936 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2968 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5936 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5935 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_742 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_2968 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2967 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2966 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2965 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVXL U5 ( .A(s3), .Z(n3) );
  CMX2X1 U6 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(s4), .Z(n2) );
endmodule


module Add_half_5937 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5938 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2969 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5938 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5937 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5939 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5940 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2970 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5940 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5939 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5941 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5942 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2971 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5942 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5941 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5943 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5944 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2972 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5944 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5943 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_743 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2972 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2971 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2970 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2969 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_5945 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_5946 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2973 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5946 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5945 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5947 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5948 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2974 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5948 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5947 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5949 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5950 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2975 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5950 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5949 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5951 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5952 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2976 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5952 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5951 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_744 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2976 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2975 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2974 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2973 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_186 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_744 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_743 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_742 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_741 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n6) );
  CIVX1 U4 ( .A(s42[0]), .Z(n4) );
  CMX2XL U5 ( .A0(s43[1]), .A1(s44[1]), .S(n6), .Z(sum4[3]) );
  CMX2XL U6 ( .A0(s43[0]), .A1(s44[0]), .S(n6), .Z(sum4[2]) );
  CMX2X1 U7 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U8 ( .A(c_out410), .Z(n3) );
  CIVX2 U9 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out4) );
  CIVX2 U12 ( .A(s41[0]), .Z(n5) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
endmodule


module Add_half_5953 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5954 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2977 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5954 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5953 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5955 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5956 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2978 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5956 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5955 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5957 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5958 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2979 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5958 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5957 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5959 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5960 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2980 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5960 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5959 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_745 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2980 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2979 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2978 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2977 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CIVX2 U7 ( .A(s1), .Z(n3) );
  CIVX2 U8 ( .A(s2), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_5961 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5962 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2981 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5962 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5961 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5963 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5964 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2982 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5964 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5963 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5965 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_5966 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2983 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5966 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5965 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5967 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5968 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2984 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5968 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5967 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_746 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_2984 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2983 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2982 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2981 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_5969 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_5970 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2985 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5970 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5969 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5971 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5972 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2986 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5972 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5971 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5973 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5974 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2987 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5974 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5973 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5975 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_5976 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENX1 U1 ( .A(n1), .B(b), .Z(sum) );
  CIVX1 U2 ( .A(a), .Z(n1) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2988 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5976 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5975 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_747 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_2988 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2987 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2986 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2985 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n6) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_5977 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5978 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2989 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5978 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5977 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5979 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5980 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2990 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5980 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5979 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5981 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_5982 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2991 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_5982 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5981 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5983 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5984 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2992 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5984 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5983 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_748 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_2992 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2991 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2990 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2989 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n4), .A1(n5), .S(n1), .Z(sum2[1]) );
  CMXI2X1 U4 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
endmodule


module bit4_187 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_748 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_747 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_746 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_745 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n6), .A1(n5), .S(n4), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
  CIVX2 U12 ( .A(s43[1]), .Z(n6) );
  CIVX2 U13 ( .A(s44[1]), .Z(n5) );
endmodule


module Add_half_5985 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5986 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2993 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5986 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5985 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5987 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5988 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2994 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5988 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5987 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5989 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5990 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2995 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5990 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5989 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5991 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5992 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2996 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5992 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5991 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_749 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_2996 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2995 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2994 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2993 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U7 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_5993 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_5994 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2997 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5994 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5993 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5995 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_5996 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_2998 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_5996 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5995 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_5997 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_5998 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_2999 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_5998 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5997 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_5999 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6000 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3000 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6000 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_5999 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_750 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_3000 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_2999 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_2998 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_2997 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_6001 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_6002 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3001 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6002 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6001 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6003 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6004 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3002 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6004 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6003 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6005 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6006 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3003 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6006 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6005 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_6007 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6008 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3004 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6008 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6007 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_751 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3004 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3003 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3002 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3001 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_6009 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(a), .B(n2), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_6010 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3005 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6010 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6009 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6011 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6012 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3006 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6012 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6011 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6013 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6014 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3007 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6014 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6013 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6015 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6016 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3008 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6016 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6015 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_752 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3008 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3007 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3006 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3005 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_188 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_752 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_751 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_750 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_749 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX1 U4 ( .A(s42[0]), .Z(n4) );
  CIVX1 U5 ( .A(s41[0]), .Z(n5) );
  CMX2XL U6 ( .A0(s43[1]), .A1(s44[1]), .S(n8), .Z(sum4[3]) );
  CMX2X1 U7 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U8 ( .A(c_out410), .Z(n3) );
  CIVX2 U9 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U10 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U11 ( .A(n1), .Z(n8) );
  CMXI2X1 U12 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n7) );
  CIVX2 U15 ( .A(s44[0]), .Z(n6) );
endmodule


module bit8_47 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n7, n8,
         n9, n10, n11, n12, n13, n14;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_188 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_187 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_186 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_185 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMXI2X2 U3 ( .A0(n9), .A1(n8), .S(c_in8), .Z(sum8[0]) );
  CIVXL U4 ( .A(s84[2]), .Z(n12) );
  CIVXL U5 ( .A(s83[2]), .Z(n13) );
  CIVX1 U6 ( .A(c_in8), .Z(n3) );
  CMX2X1 U7 ( .A0(n11), .A1(n10), .S(c_in8), .Z(n5) );
  CIVXL U8 ( .A(n14), .Z(n1) );
  CIVX2 U9 ( .A(n7), .Z(n14) );
  CIVX2 U10 ( .A(n5), .Z(sum8[1]) );
  CIVXL U11 ( .A(n1), .Z(n2) );
  CIVX1 U12 ( .A(n3), .Z(n4) );
  CMX2X2 U13 ( .A0(s81[2]), .A1(s82[2]), .S(n4), .Z(sum8[2]) );
  CMXI2XL U14 ( .A0(n13), .A1(n12), .S(n14), .Z(sum8[6]) );
  CMX2X2 U15 ( .A0(c_out810), .A1(c_out811), .S(n14), .Z(c_out8) );
  CMX2X2 U16 ( .A0(s83[0]), .A1(s84[0]), .S(n14), .Z(sum8[4]) );
  CMX2X1 U17 ( .A0(s83[3]), .A1(s84[3]), .S(n2), .Z(sum8[7]) );
  CMX2X1 U18 ( .A0(s81[3]), .A1(s82[3]), .S(n4), .Z(sum8[3]) );
  CIVXL U19 ( .A(s82[1]), .Z(n10) );
  CMX2X1 U20 ( .A0(s83[1]), .A1(s84[1]), .S(n14), .Z(sum8[5]) );
  CMXI2X1 U21 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n7) );
  CIVX2 U22 ( .A(s81[0]), .Z(n9) );
  CIVX2 U23 ( .A(s82[0]), .Z(n8) );
  CIVX2 U24 ( .A(s81[1]), .Z(n11) );
endmodule


module Add_half_6017 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_6018 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3009 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6018 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6017 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6019 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6020 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3010 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6020 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6019 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6021 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6022 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3011 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6022 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6021 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6023 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6024 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3012 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6024 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6023 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w2), .Z(n1) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_753 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3012 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3011 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3010 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3009 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s1), .Z(n5) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n6) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_6025 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6026 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3013 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6026 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6025 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_6027 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6028 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3014 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6028 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6027 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6029 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6030 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3015 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6030 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6029 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6031 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_6032 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3016 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6032 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6031 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_754 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3016 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3015 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3014 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3013 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
  CIVX2 U8 ( .A(s3), .Z(n4) );
  CIVX2 U9 ( .A(s4), .Z(n3) );
endmodule


module Add_half_6033 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6034 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3017 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6034 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6033 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6035 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6036 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3018 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6036 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6035 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6037 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6038 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3019 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6038 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6037 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6039 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6040 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3020 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6040 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6039 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_755 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3020 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3019 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3018 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3017 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6041 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6042 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3021 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6042 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6041 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6043 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6044 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3022 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6044 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6043 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6045 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6046 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3023 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6046 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6045 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6047 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6048 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3024 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6048 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6047 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_756 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3024 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3023 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3022 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3021 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_189 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_756 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_755 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_754 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_753 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n2), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n2), .Z(sum4[0]) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMX2X1 U4 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(c_out410), .A1(c_out411), .S(n1), .Z(c_out4) );
  CMX2X1 U6 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CIVX2 U7 ( .A(c_in4), .Z(n2) );
endmodule


module Add_half_6049 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_6050 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3025 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6050 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6049 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6051 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6052 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3026 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6052 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6051 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6053 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6054 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3027 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6054 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6053 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_6055 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6056 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3028 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6056 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6055 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_757 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_3028 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3027 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3026 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3025 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_6057 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_6058 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3029 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6058 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6057 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6059 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6060 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3030 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6060 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6059 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6061 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6062 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3031 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6062 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6061 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_6063 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6064 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3032 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6064 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6063 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_758 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_3032 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3031 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3030 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3029 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CIVX1 U4 ( .A(n2), .Z(n3) );
  CMXI2X1 U5 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CMX2XL U6 ( .A0(s3), .A1(s4), .S(n3), .Z(sum2[1]) );
  CMX2X1 U7 ( .A0(c_out10), .A1(c_out11), .S(n3), .Z(c_out2) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_6065 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6066 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3033 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6066 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6065 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6067 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6068 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3034 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6068 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6067 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6069 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6070 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3035 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6070 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6069 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6071 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6072 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3036 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6072 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6071 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_759 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3036 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3035 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3034 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3033 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6073 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6074 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3037 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6074 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6073 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6075 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6076 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3038 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6076 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6075 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6077 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6078 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3039 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6078 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6077 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6079 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6080 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3040 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6080 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6079 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_760 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3040 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3039 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3038 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3037 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_190 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_760 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_759 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_758 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_757 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n6), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n6), .Z(sum4[0]) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX1 U4 ( .A(c_out411), .Z(n2) );
  CIVX1 U5 ( .A(c_out410), .Z(n3) );
  CMX2X1 U6 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out4) );
  CIVX2 U10 ( .A(s43[0]), .Z(n5) );
  CIVX2 U11 ( .A(s44[0]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(n1), .Z(sum4[2]) );
  CIVX2 U13 ( .A(c_in4), .Z(n6) );
endmodule


module Add_half_6081 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6082 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3041 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6082 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6081 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6083 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6084 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3042 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6084 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6083 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6085 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6086 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3043 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6086 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6085 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6087 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6088 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3044 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6088 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6087 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_761 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3044 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3043 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3042 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3041 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6089 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6090 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3045 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6090 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6089 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6091 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6092 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3046 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6092 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6091 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6093 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6094 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3047 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6094 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6093 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6095 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6096 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3048 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6096 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6095 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_762 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3048 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3047 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3046 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3045 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6097 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6098 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3049 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6098 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6097 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6099 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6100 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3050 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6100 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6099 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6101 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6102 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3051 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6102 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6101 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6103 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6104 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3052 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6104 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6103 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_763 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3052 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3051 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3050 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3049 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6105 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6106 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3053 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6106 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6105 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6107 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6108 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3054 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6108 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6107 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6109 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6110 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3055 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6110 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6109 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6111 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6112 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3056 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6112 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6111 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_764 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3056 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3055 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3054 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3053 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_191 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_764 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_763 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_762 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_761 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_6113 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6114 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3057 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6114 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6113 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6115 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6116 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3058 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6116 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6115 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6117 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6118 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3059 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6118 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6117 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6119 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6120 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3060 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6120 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6119 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_765 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3060 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3059 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3058 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3057 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6121 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6122 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3061 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6122 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6121 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6123 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6124 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3062 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6124 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6123 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6125 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6126 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3063 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6126 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6125 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6127 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6128 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3064 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6128 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6127 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_766 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3064 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3063 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3062 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3061 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6129 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6130 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3065 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6130 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6129 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6131 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6132 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3066 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6132 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6131 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6133 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6134 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3067 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6134 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6133 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6135 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6136 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3068 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6136 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6135 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_767 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3068 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3067 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3066 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3065 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6137 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6138 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3069 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6138 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6137 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6139 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6140 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3070 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6140 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6139 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6141 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6142 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3071 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6142 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6141 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6143 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6144 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3072 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6144 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6143 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_768 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3072 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3071 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3070 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3069 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_192 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_768 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_767 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_766 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_765 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_48 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   n12, c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n5, n6, n7,
         n8, n9, n10, n11;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_192 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_191 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_190 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_189 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CAOR2X1 U8 ( .A(s84[1]), .B(n11), .C(s83[1]), .D(n9), .Z(sum8[5]) );
  CAOR2X1 U9 ( .A(s84[0]), .B(n11), .C(s83[0]), .D(n9), .Z(sum8[4]) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n10), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n10), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n10), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n10), .Z(sum8[0]) );
  CND2X1 U3 ( .A(c_out810), .B(n9), .Z(n1) );
  CND2X2 U4 ( .A(c_out811), .B(n11), .Z(n2) );
  CND2X2 U5 ( .A(n1), .B(n2), .Z(c_out8) );
  CMXI2X2 U6 ( .A0(n6), .A1(n5), .S(n11), .Z(sum8[6]) );
  CIVX1 U7 ( .A(n12), .Z(n3) );
  CIVX4 U14 ( .A(n3), .Z(sum8[7]) );
  CMXI2X1 U15 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n9) );
  CIVX2 U16 ( .A(n9), .Z(n11) );
  CIVX2 U17 ( .A(s83[2]), .Z(n6) );
  CIVX2 U18 ( .A(s84[2]), .Z(n5) );
  CIVX2 U19 ( .A(s83[3]), .Z(n8) );
  CIVX2 U20 ( .A(s84[3]), .Z(n7) );
  CMXI2X1 U21 ( .A0(n8), .A1(n7), .S(n11), .Z(n12) );
  CIVX2 U22 ( .A(c_in8), .Z(n10) );
endmodule


module bit32_12 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   n2, c1, c2, c3;

  bit8_48 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8(a32[7:0]), .b8(b32[7:0]), 
        .c_in8(c_in32) );
  bit8_47 A322 ( .sum8({sum32[15], n2, sum32[13:8]}), .c_out8(c2), .a8(
        a32[15:8]), .b8(b32[15:8]), .c_in8(c1) );
  bit8_46 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8(a32[23:16]), .b8(
        b32[23:16]), .c_in8(c2) );
  bit8_45 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8(a32[31:24]), .b8(
        b32[31:24]), .c_in8(c3) );
  CNIVX3 U1 ( .A(n2), .Z(sum32[14]) );
endmodule


module Add_half_6145 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6146 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3073 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6146 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6145 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6147 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6148 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3074 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6148 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6147 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6149 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6150 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3075 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6150 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6149 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6151 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6152 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3076 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6152 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6151 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_769 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3076 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3075 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3074 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3073 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6153 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6154 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3077 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6154 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6153 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6155 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6156 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3078 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6156 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6155 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6157 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6158 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3079 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6158 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6157 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6159 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6160 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3080 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6160 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6159 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_770 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3080 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3079 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3078 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3077 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6161 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6162 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3081 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6162 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6161 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6163 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6164 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3082 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6164 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6163 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6165 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6166 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3083 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6166 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6165 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6167 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6168 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3084 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6168 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6167 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_771 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3084 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3083 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3082 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3081 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6169 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6170 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3085 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6170 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6169 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6171 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6172 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3086 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6172 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6171 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6173 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6174 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3087 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6174 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6173 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6175 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6176 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3088 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6176 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6175 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_772 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3088 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3087 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3086 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3085 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_193 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_772 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_771 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_770 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_769 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_6177 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6178 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3089 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6178 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6177 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6179 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6180 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3090 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6180 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6179 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6181 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6182 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3091 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6182 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6181 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6183 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6184 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3092 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6184 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6183 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_773 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3092 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3091 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3090 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3089 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6185 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6186 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3093 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6186 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6185 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6187 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6188 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3094 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6188 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6187 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6189 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6190 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3095 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6190 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6189 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6191 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6192 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3096 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6192 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6191 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_774 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3096 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3095 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3094 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3093 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6193 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6194 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3097 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6194 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6193 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6195 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6196 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3098 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6196 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6195 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6197 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6198 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3099 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6198 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6197 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6199 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6200 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3100 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6200 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6199 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_775 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3100 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3099 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3098 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3097 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6201 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6202 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3101 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6202 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6201 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6203 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6204 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3102 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6204 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6203 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6205 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6206 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3103 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6206 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6205 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6207 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6208 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3104 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6208 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6207 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_776 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3104 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3103 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3102 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3101 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_194 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_776 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_775 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_774 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_773 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_6209 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6210 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3105 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6210 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6209 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6211 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6212 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3106 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6212 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6211 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6213 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6214 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3107 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6214 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6213 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6215 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6216 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3108 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6216 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6215 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_777 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3108 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3107 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3106 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3105 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6217 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6218 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3109 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6218 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6217 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6219 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6220 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3110 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6220 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6219 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6221 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6222 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3111 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6222 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6221 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6223 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6224 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3112 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6224 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6223 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_778 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3112 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3111 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3110 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3109 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6225 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6226 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3113 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6226 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6225 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6227 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6228 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3114 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6228 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6227 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6229 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6230 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3115 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6230 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6229 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6231 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6232 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3116 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6232 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6231 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_779 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3116 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3115 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3114 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3113 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6233 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6234 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3117 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6234 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6233 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6235 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6236 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3118 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6236 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6235 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6237 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6238 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3119 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6238 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6237 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6239 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6240 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3120 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6240 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6239 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_780 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3120 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3119 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3118 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3117 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_195 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_780 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_779 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_778 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_777 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_6241 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6242 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3121 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6242 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6241 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6243 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6244 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3122 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6244 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6243 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6245 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6246 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3123 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6246 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6245 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6247 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6248 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3124 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6248 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6247 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_781 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3124 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3123 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3122 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3121 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6249 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6250 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3125 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6250 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6249 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6251 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6252 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3126 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6252 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6251 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6253 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6254 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3127 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6254 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6253 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6255 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6256 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3128 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6256 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6255 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_782 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3128 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3127 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3126 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3125 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6257 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6258 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3129 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6258 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6257 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6259 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6260 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3130 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6260 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6259 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6261 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6262 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3131 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6262 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6261 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6263 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6264 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3132 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6264 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6263 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_783 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3132 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3131 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3130 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3129 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6265 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6266 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3133 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6266 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6265 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6267 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6268 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3134 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6268 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6267 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6269 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6270 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3135 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6270 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6269 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6271 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6272 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3136 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6272 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6271 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_784 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3136 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3135 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3134 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3133 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_196 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_784 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_783 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_782 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_781 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_49 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n6, n7, n8;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_196 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_195 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_194 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_193 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X4 U3 ( .A0(s83[0]), .A1(s84[0]), .S(n6), .Z(sum8[4]) );
  CMXI2XL U4 ( .A0(n8), .A1(n7), .S(n6), .Z(c_out8) );
  CMX2X2 U5 ( .A0(s81[1]), .A1(s82[1]), .S(n4), .Z(sum8[1]) );
  CMX2X1 U6 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n6) );
  CND2X2 U7 ( .A(s81[0]), .B(n1), .Z(n2) );
  CND2X1 U8 ( .A(s82[0]), .B(c_in8), .Z(n3) );
  CND2X2 U9 ( .A(n2), .B(n3), .Z(sum8[0]) );
  CIVX1 U10 ( .A(c_in8), .Z(n1) );
  CMX2X2 U11 ( .A0(s83[1]), .A1(s84[1]), .S(n6), .Z(sum8[5]) );
  CIVX2 U12 ( .A(n1), .Z(n4) );
  CMX2X1 U13 ( .A0(s81[3]), .A1(s82[3]), .S(n4), .Z(sum8[3]) );
  CMX2X1 U14 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2XL U15 ( .A0(s83[3]), .A1(s84[3]), .S(n6), .Z(sum8[7]) );
  CMX2X1 U16 ( .A0(s83[2]), .A1(s84[2]), .S(n6), .Z(sum8[6]) );
  CIVX2 U17 ( .A(c_out810), .Z(n8) );
  CIVX2 U18 ( .A(c_out811), .Z(n7) );
endmodule


module Add_half_6273 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6274 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3137 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6274 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6273 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6275 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6276 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3138 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6276 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6275 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6277 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6278 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3139 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6278 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6277 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6279 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6280 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3140 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6280 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6279 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_785 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3140 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3139 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3138 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3137 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6281 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6282 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3141 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6282 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6281 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6283 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6284 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3142 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6284 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6283 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6285 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6286 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3143 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6286 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6285 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6287 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6288 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3144 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6288 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6287 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_786 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3144 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3143 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3142 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3141 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6289 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6290 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3145 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6290 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6289 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6291 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6292 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3146 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6292 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6291 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6293 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6294 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3147 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6294 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6293 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6295 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6296 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3148 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6296 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6295 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_787 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_3148 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3147 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3146 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3145 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_6297 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6298 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3149 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6298 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6297 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6299 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6300 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3150 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6300 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6299 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6301 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6302 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3151 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6302 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6301 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_6303 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6304 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3152 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6304 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6303 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_788 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_3152 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3151 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3150 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3149 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module bit4_197 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_788 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_787 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_786 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_785 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n5), .Z(sum4[0]) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
  CIVX2 U12 ( .A(c_in4), .Z(n5) );
endmodule


module Add_half_6305 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6306 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3153 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6306 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6305 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6307 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6308 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3154 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6308 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6307 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6309 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6310 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3155 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6310 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6309 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6311 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6312 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3156 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6312 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6311 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_789 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3156 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3155 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3154 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3153 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6313 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6314 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3157 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6314 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6313 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6315 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6316 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3158 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6316 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6315 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6317 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6318 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3159 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6318 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6317 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6319 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6320 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3160 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6320 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6319 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_790 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3160 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3159 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3158 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3157 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6321 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6322 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3161 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6322 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6321 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6323 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6324 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3162 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6324 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6323 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6325 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6326 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3163 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6326 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6325 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_6327 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6328 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3164 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6328 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6327 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_791 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_3164 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3163 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3162 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3161 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMXI2X1 U3 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n4) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_6329 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6330 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3165 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6330 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6329 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6331 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6332 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3166 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6332 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6331 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6333 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6334 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3167 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6334 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6333 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_6335 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_6336 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3168 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6336 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6335 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_792 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_3168 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3167 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3166 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3165 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n5), .Z(sum2[0]) );
  CMXI2X1 U3 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n4) );
  CIVX2 U10 ( .A(c_in2), .Z(n5) );
endmodule


module bit4_198 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_792 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_791 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_790 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_789 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n11), .Z(sum4[0]) );
  CIVX2 U3 ( .A(c_out410), .Z(n3) );
  CIVX2 U4 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n8) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U8 ( .A(s41[1]), .Z(n5) );
  CIVX2 U10 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(s43[0]), .Z(n7) );
  CIVX2 U13 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX2 U15 ( .A(s43[1]), .Z(n10) );
  CIVX2 U16 ( .A(s44[1]), .Z(n9) );
  CMXI2X1 U17 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
  CIVX2 U18 ( .A(c_in4), .Z(n11) );
endmodule


module Add_half_6337 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6338 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3169 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6338 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6337 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6339 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6340 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3170 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6340 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6339 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6341 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6342 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3171 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6342 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6341 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6343 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6344 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3172 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6344 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6343 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_793 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3172 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3171 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3170 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3169 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module Add_half_6345 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6346 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3173 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6346 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6345 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6347 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6348 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3174 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6348 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6347 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6349 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6350 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3175 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6350 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6349 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6351 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6352 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3176 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6352 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6351 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_794 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3176 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3175 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3174 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3173 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U8 ( .A(s3), .Z(n5) );
  CIVX2 U9 ( .A(s4), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module Add_half_6353 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6354 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3177 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6354 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6353 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6355 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6356 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3178 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6356 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6355 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6357 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6358 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3179 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6358 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6357 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6359 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6360 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3180 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6360 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6359 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_795 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_3180 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3179 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3178 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3177 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_6361 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6362 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3181 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6362 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6361 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6363 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6364 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3182 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6364 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6363 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6365 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6366 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3183 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6366 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6365 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6367 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6368 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3184 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6368 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6367 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_796 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3184 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3183 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3182 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3181 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s3), .Z(n6) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module bit4_199 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_796 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_795 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_794 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_793 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2X1 U4 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U6 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module Add_half_6369 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6370 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3185 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6370 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6369 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6371 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6372 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3186 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6372 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6371 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6373 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6374 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3187 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6374 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6373 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6375 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6376 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3188 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6376 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6375 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_797 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3188 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3187 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3186 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3185 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(c_in2), .Z(n4) );
endmodule


module Add_half_6377 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6378 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3189 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6378 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6377 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6379 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6380 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3190 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6380 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6379 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6381 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6382 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3191 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6382 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6381 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6383 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6384 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3192 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6384 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6383 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_798 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3192 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3191 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3190 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3189 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(c_in2), .Z(n4) );
endmodule


module Add_half_6385 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6386 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3193 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6386 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6385 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6387 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6388 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3194 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6388 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6387 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6389 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6390 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3195 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6390 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6389 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6391 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6392 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3196 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6392 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6391 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_799 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3196 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3195 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3194 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3193 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_6393 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6394 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3197 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6394 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6393 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6395 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6396 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3198 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6396 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6395 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6397 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6398 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3199 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6398 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6397 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_6399 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6400 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3200 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6400 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6399 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(c_out) );
endmodule


module bit2_800 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3200 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3199 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3198 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3197 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_200 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_800 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_799 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_798 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_797 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n10), .Z(c_out4) );
  CIVX2 U4 ( .A(c_out410), .Z(n3) );
  CIVX2 U5 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n10) );
  CIVX2 U8 ( .A(s41[0]), .Z(n5) );
  CIVX2 U9 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U11 ( .A(s41[1]), .Z(n7) );
  CIVX2 U12 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U13 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n9) );
  CIVX2 U15 ( .A(s44[0]), .Z(n8) );
  CMXI2X1 U16 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CIVX2 U17 ( .A(s43[1]), .Z(n12) );
  CIVX2 U18 ( .A(s44[1]), .Z(n11) );
  CMXI2X1 U19 ( .A0(n12), .A1(n11), .S(n10), .Z(sum4[3]) );
endmodule


module bit8_50 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_200 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_199 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_198 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_197 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X1 U3 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CMX2X1 U4 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n2) );
  CIVXL U5 ( .A(s82[0]), .Z(n3) );
  CMX2X2 U6 ( .A0(s83[1]), .A1(s84[1]), .S(n2), .Z(sum8[5]) );
  CMXI2X1 U7 ( .A0(n12), .A1(n11), .S(n1), .Z(sum8[4]) );
  CMX2X2 U8 ( .A0(s83[2]), .A1(s84[2]), .S(n2), .Z(sum8[6]) );
  CMX2X1 U9 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2X1 U10 ( .A0(c_out810), .A1(c_out811), .S(n1), .Z(c_out8) );
  CMXI2X2 U11 ( .A0(n10), .A1(n9), .S(c_in8), .Z(sum8[3]) );
  CMXI2X2 U12 ( .A0(n14), .A1(n13), .S(n2), .Z(sum8[7]) );
  CND2IXL U13 ( .B(n3), .A(c_in8), .Z(n6) );
  CND2X2 U14 ( .A(n5), .B(n6), .Z(sum8[0]) );
  CIVXL U15 ( .A(c_in8), .Z(n4) );
  CND2X1 U16 ( .A(s81[0]), .B(n4), .Z(n5) );
  CMXI2X2 U17 ( .A0(n8), .A1(n7), .S(c_in8), .Z(sum8[2]) );
  CIVX2 U18 ( .A(s81[2]), .Z(n8) );
  CIVX2 U19 ( .A(s82[2]), .Z(n7) );
  CIVX2 U20 ( .A(s81[3]), .Z(n10) );
  CIVX2 U21 ( .A(s82[3]), .Z(n9) );
  CIVX2 U22 ( .A(s83[0]), .Z(n12) );
  CIVX2 U23 ( .A(s84[0]), .Z(n11) );
  CIVX2 U24 ( .A(s83[3]), .Z(n14) );
  CIVX2 U25 ( .A(s84[3]), .Z(n13) );
endmodule


module Add_half_6401 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6402 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3201 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6402 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6401 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6403 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6404 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3202 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6404 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6403 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6405 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6406 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3203 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6406 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6405 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6407 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6408 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3204 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6408 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6407 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_801 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_3204 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3203 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3202 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3201 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_6409 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6410 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3205 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6410 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6409 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6411 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6412 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3206 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6412 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6411 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6413 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6414 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3207 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6414 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6413 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6415 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6416 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3208 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6416 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6415 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_802 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_3208 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3207 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3206 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3205 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U5 ( .A(c_out10), .Z(n3) );
  CIVXL U6 ( .A(s3), .Z(n5) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
endmodule


module Add_half_6417 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6418 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3209 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6418 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6417 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6419 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6420 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3210 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6420 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6419 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6421 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6422 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3211 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6422 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6421 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6423 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6424 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3212 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6424 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6423 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_803 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_3212 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3211 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3210 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3209 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_6425 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6426 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3213 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6426 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6425 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6427 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6428 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3214 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6428 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6427 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6429 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6430 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CENXL U1 ( .A(a), .B(b), .Z(n1) );
  CIVX1 U2 ( .A(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3215 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6430 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6429 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6431 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6432 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3216 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6432 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6431 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_804 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3216 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3215 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3214 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3213 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_201 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_804 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_803 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_802 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_801 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(c_out410), .A1(c_out411), .S(n2), .Z(c_out4) );
  CMX2XL U4 ( .A0(s43[1]), .A1(s44[1]), .S(n2), .Z(sum4[3]) );
  CMX2XL U5 ( .A0(s43[0]), .A1(s44[0]), .S(n2), .Z(sum4[2]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U7 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n2) );
endmodule


module Add_half_6433 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6434 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3217 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6434 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6433 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6435 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6436 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3218 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6436 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6435 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6437 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6438 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3219 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6438 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6437 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6439 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6440 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3220 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6440 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6439 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_805 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_3220 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3219 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3218 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3217 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
endmodule


module Add_half_6441 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6442 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3221 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6442 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6441 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6443 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6444 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3222 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6444 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6443 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6445 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6446 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3223 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6446 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6445 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6447 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6448 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3224 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6448 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6447 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_806 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_3224 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3223 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3222 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3221 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
endmodule


module Add_half_6449 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6450 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3225 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6450 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6449 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6451 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6452 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3226 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6452 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6451 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6453 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6454 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3227 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6454 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6453 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6455 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6456 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3228 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6456 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6455 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_807 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3228 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3227 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3226 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3225 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_6457 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6458 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3229 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6458 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6457 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6459 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6460 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3230 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6460 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6459 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6461 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6462 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3231 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6462 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6461 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6463 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6464 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3232 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6464 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6463 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_808 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3232 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3231 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3230 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3229 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_202 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_808 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_807 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_806 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_805 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n3), .A1(n2), .S(n10), .Z(c_out4) );
  CIVX2 U4 ( .A(c_out410), .Z(n3) );
  CIVX2 U5 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n10) );
  CIVX2 U8 ( .A(s41[0]), .Z(n5) );
  CIVX2 U9 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U11 ( .A(s41[1]), .Z(n7) );
  CIVX2 U12 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U13 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n9) );
  CIVX2 U15 ( .A(s44[0]), .Z(n8) );
  CMXI2X1 U16 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CIVX2 U17 ( .A(s43[1]), .Z(n12) );
  CIVX2 U18 ( .A(s44[1]), .Z(n11) );
  CMXI2X1 U19 ( .A0(n12), .A1(n11), .S(n10), .Z(sum4[3]) );
endmodule


module Add_half_6465 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6466 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3233 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6466 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6465 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6467 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6468 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3234 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6468 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6467 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6469 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6470 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3235 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6470 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6469 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6471 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6472 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3236 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6472 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6471 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_809 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3236 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3235 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3234 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3233 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n2) );
  CIVX2 U7 ( .A(s3), .Z(n4) );
  CIVX2 U8 ( .A(s4), .Z(n3) );
  CMXI2X1 U9 ( .A0(n4), .A1(n3), .S(n2), .Z(sum2[1]) );
endmodule


module Add_half_6473 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6474 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3237 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6474 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6473 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6475 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6476 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3238 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6476 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6475 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6477 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6478 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3239 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6478 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6477 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6479 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6480 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3240 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6480 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6479 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_810 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_3240 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3239 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3238 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3237 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_6481 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6482 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3241 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6482 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6481 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6483 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6484 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3242 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6484 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6483 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6485 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6486 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3243 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6486 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6485 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6487 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6488 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3244 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6488 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6487 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_811 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3244 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3243 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3242 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3241 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_6489 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_6490 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3245 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6490 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6489 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6491 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6492 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3246 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6492 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6491 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6493 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6494 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3247 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6494 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6493 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6495 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6496 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3248 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6496 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6495 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_812 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3248 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3247 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3246 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3245 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_203 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_812 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_811 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_810 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_809 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out4) );
  CIVX1 U4 ( .A(s42[0]), .Z(n4) );
  CMX2XL U5 ( .A0(s43[1]), .A1(s44[1]), .S(n8), .Z(sum4[3]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n8) );
  CIVX2 U11 ( .A(s41[0]), .Z(n5) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U13 ( .A(s43[0]), .Z(n7) );
  CIVX2 U14 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U15 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
endmodule


module Add_half_6497 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6498 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3249 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6498 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6497 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6499 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6500 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3250 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6500 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6499 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6501 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6502 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3251 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6502 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6501 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6503 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6504 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3252 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6504 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6503 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_813 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3252 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3251 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3250 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3249 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CIVX2 U7 ( .A(s1), .Z(n3) );
  CIVX2 U8 ( .A(s2), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_6505 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6506 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3253 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6506 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6505 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6507 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6508 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3254 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6508 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6507 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6509 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_6510 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3255 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6510 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6509 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6511 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6512 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3256 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6512 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6511 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_814 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_3256 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3255 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3254 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3253 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_6513 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6514 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3257 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6514 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6513 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6515 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6516 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3258 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6516 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6515 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6517 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6518 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3259 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6518 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6517 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6519 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6520 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3260 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6520 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6519 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_815 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3260 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3259 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3258 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3257 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_6521 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6522 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3261 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6522 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6521 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6523 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6524 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3262 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6524 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6523 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6525 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_6526 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3263 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6526 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6525 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX1 U1 ( .A(w3), .Z(n2) );
  CND2X1 U2 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6527 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6528 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3264 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6528 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6527 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_816 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3264 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3263 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3262 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3261 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_204 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_816 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_815 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_814 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_813 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2X1 U3 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out4) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n6), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CIVX2 U7 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n6) );
  CIVX2 U10 ( .A(s41[1]), .Z(n5) );
  CIVX2 U11 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U12 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U13 ( .A(s43[1]), .Z(n8) );
  CIVX2 U14 ( .A(s44[1]), .Z(n7) );
  CMXI2X1 U15 ( .A0(n8), .A1(n7), .S(n6), .Z(sum4[3]) );
endmodule


module bit8_51 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_204 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_203 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_202 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_201 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CND2X4 U3 ( .A(n3), .B(n4), .Z(c_out8) );
  CIVX1 U4 ( .A(n7), .Z(n12) );
  CMX2X1 U5 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n1) );
  CMX2X2 U6 ( .A0(s81[3]), .A1(s82[3]), .S(n6), .Z(sum8[3]) );
  CMX2X2 U7 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CIVXL U8 ( .A(c_in8), .Z(n5) );
  CND2X2 U9 ( .A(n2), .B(c_out810), .Z(n3) );
  CND2X1 U10 ( .A(c_out811), .B(n12), .Z(n4) );
  CIVX1 U11 ( .A(n12), .Z(n2) );
  CMX2X2 U12 ( .A0(s83[1]), .A1(s84[1]), .S(n1), .Z(sum8[5]) );
  CMX2X2 U13 ( .A0(s83[2]), .A1(s84[2]), .S(n1), .Z(sum8[6]) );
  CIVXL U14 ( .A(n5), .Z(n6) );
  CMXI2X1 U15 ( .A0(n9), .A1(n8), .S(c_in8), .Z(sum8[0]) );
  CMXI2X1 U16 ( .A0(n11), .A1(n10), .S(n12), .Z(sum8[4]) );
  CMX2X1 U17 ( .A0(s83[3]), .A1(s84[3]), .S(n1), .Z(sum8[7]) );
  CMX2X1 U18 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMXI2X1 U19 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n7) );
  CIVX2 U20 ( .A(s81[0]), .Z(n9) );
  CIVX2 U21 ( .A(s82[0]), .Z(n8) );
  CIVX2 U22 ( .A(s83[0]), .Z(n11) );
  CIVX2 U23 ( .A(s84[0]), .Z(n10) );
endmodule


module Add_half_6529 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6530 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3265 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6530 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6529 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6531 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6532 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3266 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6532 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6531 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6533 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6534 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3267 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6534 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6533 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6535 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6536 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3268 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6536 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6535 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_817 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_3268 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3267 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3266 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3265 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_6537 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6538 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3269 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6538 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6537 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6539 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6540 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3270 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6540 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6539 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6541 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6542 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3271 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6542 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6541 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6543 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6544 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3272 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6544 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6543 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_818 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_3272 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3271 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3270 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3269 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n2) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module Add_half_6545 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6546 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3273 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6546 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6545 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6547 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX2 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6548 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3274 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6548 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6547 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6549 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6550 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3275 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6550 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6549 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX1 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6551 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6552 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3276 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6552 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6551 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_819 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_3276 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3275 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3274 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3273 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U4 ( .A(c_in2), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n3) );
  CMXI2X1 U6 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CIVX1 U7 ( .A(c_out11), .Z(n4) );
  CIVX1 U8 ( .A(c_out10), .Z(n5) );
  CMX2XL U9 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U10 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_6553 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6554 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3277 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6554 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6553 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6555 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6556 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3278 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6556 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6555 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6557 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6558 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3279 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6558 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6557 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6559 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6560 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3280 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6560 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6559 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_820 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3280 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3279 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3278 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3277 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CIVXL U4 ( .A(n1), .Z(n4) );
  CMXI2X1 U5 ( .A0(n2), .A1(n3), .S(n1), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U7 ( .A(c_out10), .Z(n3) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
endmodule


module bit4_205 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_820 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_819 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_818 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_817 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CANR2X1 U3 ( .A(c_out400), .B(n3), .C(c_in4), .D(c_out401), .Z(n2) );
  CIVX1 U4 ( .A(s42[0]), .Z(n6) );
  CNIVXL U5 ( .A(n2), .Z(n1) );
  CANR2X1 U6 ( .A(n3), .B(c_out400), .C(c_in4), .D(c_out401), .Z(n12) );
  CIVX1 U7 ( .A(c_out410), .Z(n4) );
  CIVX1 U8 ( .A(c_out411), .Z(n5) );
  CIVX1 U9 ( .A(s44[1]), .Z(n14) );
  CIVX1 U10 ( .A(s41[0]), .Z(n7) );
  CMXI2XL U11 ( .A0(n14), .A1(n13), .S(n1), .Z(sum4[3]) );
  CIVX2 U12 ( .A(c_in4), .Z(n3) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(n12), .Z(c_out4) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U15 ( .A(s41[1]), .Z(n9) );
  CIVX2 U16 ( .A(s42[1]), .Z(n8) );
  CMXI2X1 U17 ( .A0(n9), .A1(n8), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U18 ( .A(s44[0]), .Z(n11) );
  CIVX2 U19 ( .A(s43[0]), .Z(n10) );
  CMXI2X1 U20 ( .A0(n11), .A1(n10), .S(n2), .Z(sum4[2]) );
  CIVX2 U21 ( .A(s43[1]), .Z(n13) );
endmodule


module Add_half_6561 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6562 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3281 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6562 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6561 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6563 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6564 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3282 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6564 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6563 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6565 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6566 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3283 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6566 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6565 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6567 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6568 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3284 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6568 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6567 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_821 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3284 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3283 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3282 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3281 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_6569 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6570 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3285 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6570 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6569 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6571 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6572 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3286 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6572 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6571 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6573 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6574 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3287 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6574 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6573 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6575 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6576 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3288 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6576 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6575 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_822 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_3288 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3287 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3286 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3285 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2XL U4 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CIVX1 U5 ( .A(s2), .Z(n2) );
  CIVX1 U6 ( .A(s1), .Z(n3) );
  CMX2X1 U7 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
endmodule


module Add_half_6577 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_6578 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3289 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6578 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6577 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6579 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6580 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3290 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6580 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6579 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6581 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_6582 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3291 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6582 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6581 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module Add_half_6583 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6584 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3292 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6584 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6583 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_823 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_3292 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3291 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3290 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3289 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X2 U3 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n1) );
  CIVX2 U4 ( .A(c_in2), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out01), .A1(c_out00), .S(n2), .Z(n3) );
  CMX2X1 U6 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMXI2X1 U7 ( .A0(n4), .A1(n5), .S(n3), .Z(c_out2) );
  CIVX1 U8 ( .A(c_out11), .Z(n4) );
  CMX2X1 U9 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U10 ( .A(c_out10), .Z(n5) );
endmodule


module Add_half_6585 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6586 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3293 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6586 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6585 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6587 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6588 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3294 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6588 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6587 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6589 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6590 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3295 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6590 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6589 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6591 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6592 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3296 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6592 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6591 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w2), .Z(n1) );
  CIVX2 U3 ( .A(w3), .Z(n2) );
endmodule


module bit2_824 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_3296 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3295 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3294 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3293 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVXL U4 ( .A(s1), .Z(n6) );
  CMXI2X1 U5 ( .A0(n3), .A1(n4), .S(n2), .Z(c_out2) );
  CMXI2XL U6 ( .A0(n8), .A1(n7), .S(n1), .Z(sum2[1]) );
  CIVX1 U7 ( .A(c_out10), .Z(n4) );
  CIVX2 U8 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U9 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n2) );
  CIVX2 U10 ( .A(s2), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U12 ( .A(s3), .Z(n8) );
  CIVX2 U13 ( .A(s4), .Z(n7) );
endmodule


module bit4_206 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_824 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_823 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_822 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_821 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CND2X2 U3 ( .A(c_out411), .B(n1), .Z(n2) );
  CND2X1 U4 ( .A(c_out410), .B(n7), .Z(n3) );
  CND2X2 U5 ( .A(n2), .B(n3), .Z(c_out4) );
  CIVX2 U6 ( .A(n7), .Z(n1) );
  CND2X1 U7 ( .A(n5), .B(n6), .Z(sum4[2]) );
  CND2X1 U8 ( .A(n4), .B(s44[0]), .Z(n5) );
  CIVX1 U9 ( .A(n8), .Z(n4) );
  CANR2X1 U10 ( .A(c_out400), .B(n9), .C(c_in4), .D(c_out401), .Z(n8) );
  CND2XL U11 ( .A(n8), .B(s43[0]), .Z(n6) );
  CANR2X1 U12 ( .A(c_out400), .B(n9), .C(c_in4), .D(c_out401), .Z(n7) );
  CANR2XL U13 ( .A(n9), .B(c_out400), .C(c_in4), .D(c_out401), .Z(n10) );
  CMX2X1 U14 ( .A0(s44[1]), .A1(s43[1]), .S(n10), .Z(sum4[3]) );
  CMX2X1 U15 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U16 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U17 ( .A(c_in4), .Z(n9) );
endmodule


module Add_half_6593 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6594 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3297 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6594 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6593 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6595 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6596 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3298 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6596 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6595 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6597 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6598 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3299 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6598 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6597 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6599 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6600 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3300 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6600 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6599 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_825 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3300 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3299 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3298 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3297 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6601 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6602 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3301 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6602 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6601 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6603 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6604 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3302 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6604 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6603 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6605 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6606 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3303 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6606 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6605 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6607 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6608 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3304 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6608 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6607 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_826 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3304 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3303 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3302 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3301 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6609 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6610 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3305 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6610 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6609 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6611 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6612 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3306 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6612 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6611 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6613 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6614 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3307 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6614 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6613 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6615 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6616 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3308 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6616 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6615 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_827 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3308 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3307 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3306 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3305 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6617 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6618 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3309 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6618 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6617 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6619 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6620 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3310 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6620 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6619 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6621 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6622 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3311 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6622 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6621 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6623 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6624 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3312 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6624 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6623 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_828 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3312 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3311 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3310 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3309 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_207 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_828 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_827 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_826 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_825 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_6625 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6626 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3313 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6626 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6625 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6627 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6628 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3314 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6628 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6627 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6629 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6630 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3315 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6630 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6629 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6631 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6632 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3316 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6632 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6631 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_829 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3316 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3315 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3314 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3313 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6633 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6634 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3317 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6634 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6633 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6635 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6636 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3318 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6636 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6635 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6637 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6638 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3319 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6638 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6637 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6639 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6640 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3320 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6640 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6639 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_830 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3320 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3319 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3318 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3317 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6641 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6642 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3321 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6642 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6641 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6643 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6644 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3322 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6644 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6643 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6645 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6646 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3323 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6646 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6645 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6647 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6648 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3324 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6648 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6647 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_831 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3324 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3323 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3322 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3321 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6649 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6650 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3325 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6650 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6649 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6651 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6652 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3326 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6652 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6651 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6653 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6654 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3327 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6654 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6653 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6655 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6656 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3328 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6656 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6655 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_832 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3328 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3327 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3326 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3325 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_208 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_832 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_831 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_830 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_829 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_52 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8, n9;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_208 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_207 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_206 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_205 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CAOR2X1 U10 ( .A(s82[3]), .B(c_in8), .C(s81[3]), .D(n9), .Z(sum8[3]) );
  CAOR2X1 U11 ( .A(s82[2]), .B(c_in8), .C(s81[2]), .D(n9), .Z(sum8[2]) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n9), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n9), .Z(sum8[0]) );
  CIVX1 U3 ( .A(s83[2]), .Z(n7) );
  CND2X2 U4 ( .A(c_out811), .B(n8), .Z(n2) );
  CND2X4 U5 ( .A(n1), .B(n2), .Z(c_out8) );
  CND2X2 U6 ( .A(c_out810), .B(n3), .Z(n1) );
  CIVX1 U7 ( .A(s84[0]), .Z(n4) );
  CMX2X2 U8 ( .A0(s84[1]), .A1(s83[1]), .S(n3), .Z(sum8[5]) );
  CMXI2X1 U9 ( .A0(n6), .A1(n7), .S(n3), .Z(sum8[6]) );
  CIVX1 U14 ( .A(s84[2]), .Z(n6) );
  CMX2X2 U15 ( .A0(s83[3]), .A1(s84[3]), .S(n8), .Z(sum8[7]) );
  CMXI2X4 U16 ( .A0(n5), .A1(n4), .S(n8), .Z(sum8[4]) );
  CIVX1 U17 ( .A(s83[0]), .Z(n5) );
  CMXI2X1 U18 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n3) );
  CIVX2 U19 ( .A(n3), .Z(n8) );
  CIVX2 U20 ( .A(c_in8), .Z(n9) );
endmodule


module bit32_13 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   c1, c2, c3;

  bit8_52 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8(a32[7:0]), .b8(b32[7:0]), 
        .c_in8(c_in32) );
  bit8_51 A322 ( .sum8(sum32[15:8]), .c_out8(c2), .a8(a32[15:8]), .b8(
        b32[15:8]), .c_in8(c1) );
  bit8_50 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8(a32[23:16]), .b8(
        b32[23:16]), .c_in8(c2) );
  bit8_49 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8(a32[31:24]), .b8(
        b32[31:24]), .c_in8(c3) );
endmodule


module Add_half_6657 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6658 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3329 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6658 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6657 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6659 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6660 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3330 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6660 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6659 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6661 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6662 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3331 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6662 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6661 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6663 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6664 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3332 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6664 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6663 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_833 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3332 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3331 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3330 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3329 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6665 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6666 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3333 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6666 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6665 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6667 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6668 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3334 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6668 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6667 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6669 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6670 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3335 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6670 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6669 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6671 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6672 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3336 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6672 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6671 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_834 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3336 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3335 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3334 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3333 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6673 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6674 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3337 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6674 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6673 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6675 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6676 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3338 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6676 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6675 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6677 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6678 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3339 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6678 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6677 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6679 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6680 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3340 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6680 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6679 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_835 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3340 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3339 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3338 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3337 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6681 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6682 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3341 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6682 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6681 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6683 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6684 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3342 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6684 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6683 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6685 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6686 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3343 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6686 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6685 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6687 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6688 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3344 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6688 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6687 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_836 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3344 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3343 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3342 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3341 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_209 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_836 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_835 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_834 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_833 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_6689 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6690 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3345 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6690 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6689 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6691 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6692 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3346 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6692 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6691 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6693 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6694 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3347 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6694 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6693 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6695 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6696 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3348 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6696 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6695 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_837 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3348 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3347 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3346 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3345 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6697 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6698 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3349 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6698 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6697 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6699 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6700 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3350 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6700 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6699 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6701 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6702 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3351 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6702 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6701 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6703 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6704 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3352 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6704 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6703 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_838 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3352 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3351 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3350 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3349 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6705 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6706 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3353 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6706 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6705 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6707 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6708 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3354 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6708 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6707 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6709 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6710 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3355 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6710 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6709 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6711 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6712 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3356 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6712 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6711 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_839 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3356 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3355 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3354 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3353 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6713 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6714 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3357 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6714 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6713 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6715 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6716 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3358 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6716 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6715 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6717 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6718 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3359 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6718 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6717 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6719 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6720 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3360 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6720 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6719 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_840 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3360 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3359 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3358 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3357 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_210 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_840 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_839 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_838 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_837 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_6721 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6722 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3361 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6722 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6721 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6723 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6724 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3362 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6724 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6723 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6725 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6726 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3363 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6726 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6725 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6727 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6728 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3364 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6728 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6727 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_841 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3364 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3363 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3362 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3361 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6729 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6730 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3365 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6730 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6729 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6731 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6732 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3366 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6732 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6731 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6733 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6734 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3367 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6734 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6733 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6735 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6736 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3368 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6736 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6735 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_842 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3368 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3367 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3366 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3365 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6737 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6738 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3369 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6738 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6737 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6739 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6740 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3370 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6740 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6739 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6741 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6742 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3371 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6742 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6741 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6743 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6744 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3372 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6744 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6743 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_843 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3372 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3371 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3370 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3369 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6745 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6746 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3373 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6746 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6745 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6747 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6748 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3374 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6748 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6747 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6749 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6750 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3375 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6750 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6749 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6751 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6752 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3376 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6752 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6751 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_844 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3376 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3375 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3374 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3373 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_211 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_844 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_843 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_842 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_841 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_6753 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6754 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3377 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6754 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6753 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6755 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6756 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3378 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6756 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6755 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6757 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6758 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3379 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6758 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6757 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6759 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6760 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3380 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6760 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6759 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_845 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3380 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3379 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3378 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3377 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6761 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6762 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3381 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6762 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6761 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6763 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6764 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3382 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6764 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6763 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6765 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6766 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3383 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6766 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6765 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6767 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6768 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3384 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6768 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6767 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_846 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3384 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3383 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3382 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3381 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6769 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6770 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3385 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6770 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6769 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6771 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6772 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3386 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6772 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6771 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6773 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6774 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3387 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6774 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6773 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6775 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6776 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3388 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6776 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6775 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_847 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3388 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3387 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3386 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3385 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6777 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6778 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3389 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6778 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6777 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6779 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6780 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3390 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6780 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6779 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6781 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6782 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3391 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6782 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6781 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6783 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6784 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3392 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6784 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6783 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_848 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3392 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3391 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3390 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3389 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_212 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_848 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_847 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_846 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_845 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module bit8_53 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8, n9;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_212 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_211 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_210 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_209 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X2 U3 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n7) );
  CMX2X2 U4 ( .A0(s81[3]), .A1(s82[3]), .S(c_in8), .Z(sum8[3]) );
  CMX2X2 U5 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CMX2X2 U6 ( .A0(s81[0]), .A1(s82[0]), .S(c_in8), .Z(sum8[0]) );
  CND2X1 U7 ( .A(s83[3]), .B(n1), .Z(n2) );
  CND2XL U8 ( .A(s84[3]), .B(n7), .Z(n3) );
  CND2X2 U9 ( .A(n2), .B(n3), .Z(sum8[7]) );
  CIVXL U10 ( .A(n7), .Z(n1) );
  CND2X1 U11 ( .A(s81[1]), .B(n4), .Z(n5) );
  CND2XL U12 ( .A(s82[1]), .B(c_in8), .Z(n6) );
  CND2X2 U13 ( .A(n5), .B(n6), .Z(sum8[1]) );
  CIVXL U14 ( .A(c_in8), .Z(n4) );
  CMX2X2 U15 ( .A0(s83[0]), .A1(s84[0]), .S(n7), .Z(sum8[4]) );
  CMX2X1 U16 ( .A0(s83[2]), .A1(s84[2]), .S(n7), .Z(sum8[6]) );
  CMX2X1 U17 ( .A0(s83[1]), .A1(s84[1]), .S(n7), .Z(sum8[5]) );
  CMXI2XL U18 ( .A0(n9), .A1(n8), .S(n7), .Z(c_out8) );
  CIVX2 U19 ( .A(c_out810), .Z(n9) );
  CIVX2 U20 ( .A(c_out811), .Z(n8) );
endmodule


module Add_half_6785 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6786 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3393 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6786 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6785 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6787 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6788 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3394 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6788 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6787 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6789 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6790 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3395 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6790 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6789 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6791 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6792 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3396 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6792 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6791 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_849 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3396 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3395 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3394 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3393 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6793 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6794 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3397 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6794 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6793 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6795 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6796 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3398 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6796 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6795 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6797 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6798 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3399 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6798 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6797 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6799 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6800 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3400 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6800 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6799 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_850 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3400 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3399 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3398 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3397 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6801 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6802 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3401 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6802 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6801 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6803 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6804 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3402 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6804 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6803 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6805 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6806 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3403 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6806 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6805 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6807 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6808 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3404 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6808 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6807 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_851 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3404 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3403 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3402 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3401 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6809 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6810 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3405 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6810 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6809 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6811 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6812 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3406 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6812 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6811 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6813 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6814 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3407 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6814 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6813 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6815 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6816 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3408 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6816 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6815 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_852 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3408 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3407 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3406 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3405 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_213 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_852 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_851 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_850 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_849 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_6817 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6818 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3409 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6818 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6817 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6819 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6820 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3410 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6820 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6819 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6821 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6822 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3411 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6822 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6821 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6823 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6824 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3412 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6824 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6823 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_853 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3412 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3411 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3410 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3409 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6825 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6826 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3413 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6826 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6825 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6827 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6828 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3414 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6828 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6827 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6829 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6830 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3415 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6830 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6829 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6831 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6832 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3416 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6832 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6831 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_854 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3416 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3415 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3414 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3413 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6833 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6834 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3417 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6834 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6833 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6835 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6836 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3418 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6836 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6835 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6837 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6838 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3419 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6838 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6837 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6839 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6840 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3420 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6840 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6839 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_855 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3420 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3419 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3418 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3417 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_6841 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6842 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3421 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6842 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6841 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6843 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6844 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3422 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6844 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6843 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6845 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6846 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3423 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6846 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6845 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6847 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6848 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3424 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6848 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6847 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_856 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3424 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3423 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3422 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3421 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_214 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_856 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_855 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_854 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_853 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in4), .Z(n4) );
  CAOR2X1 U6 ( .A(s44[1]), .B(n5), .C(s43[1]), .D(n1), .Z(sum4[3]) );
  CAOR2X1 U7 ( .A(s44[0]), .B(n5), .C(s43[0]), .D(n1), .Z(sum4[2]) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CAOR2X1 U10 ( .A(c_out411), .B(n5), .C(c_out410), .D(n1), .Z(c_out4) );
  CANR2X1 U3 ( .A(c_out401), .B(c_in4), .C(c_out400), .D(n4), .Z(n1) );
endmodule


module Add_half_6849 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6850 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3425 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6850 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6849 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6851 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6852 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3426 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6852 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6851 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6853 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_6854 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3427 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6854 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6853 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_6855 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_6856 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3428 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6856 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6855 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_857 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_3428 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3427 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3426 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3425 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n7), .Z(sum2[0]) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX2 U12 ( .A(c_in2), .Z(n7) );
endmodule


module Add_half_6857 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6858 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3429 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6858 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6857 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6859 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6860 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3430 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6860 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6859 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6861 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_6862 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3431 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6862 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6861 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CNR2X1 U1 ( .A(w3), .B(w2), .Z(n1) );
  CIVX2 U2 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_6863 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_6864 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3432 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6864 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6863 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_858 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3432 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3431 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3430 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3429 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n6), .Z(sum2[0]) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n5) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
  CIVX2 U11 ( .A(c_in2), .Z(n6) );
endmodule


module Add_half_6865 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6866 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3433 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6866 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6865 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6867 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6868 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3434 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6868 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6867 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6869 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6870 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3435 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6870 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6869 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6871 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6872 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3436 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6872 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6871 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_859 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_3436 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3435 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3434 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3433 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_6873 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6874 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3437 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6874 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6873 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6875 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6876 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3438 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6876 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6875 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6877 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6878 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3439 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6878 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6877 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6879 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6880 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3440 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6880 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6879 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_860 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3440 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3439 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3438 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3437 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s3), .Z(n6) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module bit4_215 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_860 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_859 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_858 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_857 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2XL U4 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2X1 U5 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module Add_half_6881 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6882 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3441 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6882 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6881 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6883 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6884 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3442 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6884 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6883 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6885 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX1 U1 ( .A(n1), .Z(c_out) );
  CND2X1 U2 ( .A(a), .B(b), .Z(n1) );
  CEOXL U3 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6886 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3443 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6886 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6885 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6887 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6888 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3444 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6888 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6887 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_861 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3444 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3443 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3442 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3441 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(c_in2), .Z(n4) );
endmodule


module Add_half_6889 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6890 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3445 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6890 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6889 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6891 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_6892 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3446 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6892 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6891 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_6893 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CND2X1 U1 ( .A(a), .B(b), .Z(n1) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(n1), .Z(c_out) );
endmodule


module Add_half_6894 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3447 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6894 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6893 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6895 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6896 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(a), .Z(n1) );
  CENX1 U3 ( .A(b), .B(n1), .Z(sum) );
endmodule


module Add_full_3448 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6896 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6895 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_862 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3448 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3447 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3446 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3445 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U9 ( .A(c_in2), .Z(n4) );
endmodule


module Add_half_6897 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6898 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3449 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6898 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6897 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6899 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6900 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3450 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6900 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6899 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6901 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6902 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3451 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6902 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6901 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6903 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6904 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3452 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6904 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6903 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_863 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3452 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3451 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3450 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3449 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_6905 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6906 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3453 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6906 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6905 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6907 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6908 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3454 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6908 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6907 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6909 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6910 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3455 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6910 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6909 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6911 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6912 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3456 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6912 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6911 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_864 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3456 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3455 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3454 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3453 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_216 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_864 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_863 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_862 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_861 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX2 U3 ( .A(c_out410), .Z(n3) );
  CIVX2 U4 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n10) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n10), .Z(c_out4) );
  CIVX2 U8 ( .A(s41[0]), .Z(n5) );
  CIVX2 U9 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U11 ( .A(s41[1]), .Z(n7) );
  CIVX2 U12 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U13 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U14 ( .A(s43[0]), .Z(n9) );
  CIVX2 U15 ( .A(s44[0]), .Z(n8) );
  CMXI2X1 U16 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CIVX2 U17 ( .A(s43[1]), .Z(n12) );
  CIVX2 U18 ( .A(s44[1]), .Z(n11) );
  CMXI2X1 U19 ( .A0(n12), .A1(n11), .S(n10), .Z(sum4[3]) );
endmodule


module bit8_54 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_216 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_215 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_214 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_213 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CND2X2 U3 ( .A(c_out810), .B(n8), .Z(n9) );
  CMX2X2 U4 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n4) );
  CIVX2 U5 ( .A(n5), .Z(n1) );
  CIVX2 U6 ( .A(c_in8), .Z(n5) );
  CIVX1 U7 ( .A(s81[0]), .Z(n2) );
  CND2IX1 U8 ( .B(n2), .A(n5), .Z(n6) );
  CMX2X2 U9 ( .A0(s81[2]), .A1(s82[2]), .S(c_in8), .Z(sum8[2]) );
  CND2X1 U10 ( .A(c_out811), .B(n4), .Z(n10) );
  CIVX2 U11 ( .A(n4), .Z(n8) );
  CMX2X2 U12 ( .A0(s81[1]), .A1(s82[1]), .S(n1), .Z(sum8[1]) );
  CMXI2X1 U13 ( .A0(n13), .A1(n14), .S(n3), .Z(sum8[4]) );
  CMXI2X1 U14 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n3) );
  CMX2X2 U15 ( .A0(s84[2]), .A1(s83[2]), .S(n8), .Z(sum8[6]) );
  CND2XL U16 ( .A(c_in8), .B(s82[0]), .Z(n7) );
  CND2X2 U17 ( .A(n6), .B(n7), .Z(sum8[0]) );
  CMX2X1 U18 ( .A0(s83[3]), .A1(s84[3]), .S(n4), .Z(sum8[7]) );
  CND2X2 U19 ( .A(n9), .B(n10), .Z(c_out8) );
  CMX2X1 U20 ( .A0(s83[1]), .A1(s84[1]), .S(n4), .Z(sum8[5]) );
  CMXI2X2 U21 ( .A0(n12), .A1(n11), .S(c_in8), .Z(sum8[3]) );
  CIVX2 U22 ( .A(s81[3]), .Z(n12) );
  CIVX2 U23 ( .A(s82[3]), .Z(n11) );
  CIVX2 U24 ( .A(s83[0]), .Z(n14) );
  CIVX2 U25 ( .A(s84[0]), .Z(n13) );
endmodule


module Add_half_6913 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6914 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3457 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6914 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6913 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6915 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6916 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3458 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6916 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6915 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6917 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6918 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3459 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6918 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6917 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6919 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6920 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3460 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6920 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6919 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_865 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7;

  Add_full_3460 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3459 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3458 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3457 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n7), .A1(n6), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n7) );
  CIVX2 U12 ( .A(s4), .Z(n6) );
endmodule


module Add_half_6921 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6922 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3461 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6922 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6921 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6923 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6924 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3462 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6924 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6923 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6925 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6926 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3463 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6926 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6925 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6927 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6928 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3464 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6928 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6927 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_866 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_3464 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3463 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3462 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3461 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n5), .A1(n4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX1 U5 ( .A(c_out10), .Z(n3) );
  CIVXL U6 ( .A(s3), .Z(n5) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
  CIVX2 U10 ( .A(s4), .Z(n4) );
endmodule


module Add_half_6929 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6930 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3465 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6930 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6929 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6931 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6932 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3466 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6932 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6931 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6933 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6934 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3467 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6934 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6933 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6935 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6936 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3468 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6936 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6935 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_867 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_3468 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3467 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3466 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3465 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_6937 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6938 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3469 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6938 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6937 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6939 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6940 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3470 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6940 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6939 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6941 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6942 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3471 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6942 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6941 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6943 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6944 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3472 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6944 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6943 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_868 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3472 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3471 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3470 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3469 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_217 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_868 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_867 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_866 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_865 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n2), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n2), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(c_out410), .A1(c_out411), .S(n2), .Z(c_out4) );
  CMX2X1 U6 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U7 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CMXI2X1 U8 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U9 ( .A(n1), .Z(n2) );
endmodule


module Add_half_6945 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6946 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3473 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6946 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6945 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6947 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6948 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3474 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6948 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6947 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6949 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6950 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3475 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6950 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6949 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6951 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6952 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3476 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6952 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6951 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_869 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_3476 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3475 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3474 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3473 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
endmodule


module Add_half_6953 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6954 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3477 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6954 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6953 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6955 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_6956 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3478 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6956 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6955 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6957 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6958 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3479 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_6958 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6957 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6959 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6960 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3480 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6960 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6959 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_870 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_3480 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3479 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3478 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3477 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out2) );
endmodule


module Add_half_6961 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6962 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3481 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6962 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6961 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6963 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6964 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3482 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6964 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6963 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6965 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6966 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3483 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6966 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6965 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_6967 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6968 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3484 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_6968 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6967 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_871 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3484 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3483 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3482 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3481 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n6) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_6969 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6970 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3485 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6970 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6969 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6971 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6972 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3486 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6972 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6971 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6973 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6974 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3487 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6974 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6973 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6975 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6976 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3488 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6976 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6975 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_872 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3488 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3487 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3486 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3485 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_218 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_872 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_871 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_870 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_869 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U4 ( .A(c_out410), .Z(n3) );
  CIVX2 U5 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n8) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n8), .Z(c_out4) );
  CIVX2 U9 ( .A(s41[1]), .Z(n5) );
  CIVX2 U10 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U12 ( .A(s43[0]), .Z(n7) );
  CIVX2 U13 ( .A(s44[0]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n8), .Z(sum4[2]) );
  CIVX2 U15 ( .A(s43[1]), .Z(n10) );
  CIVX2 U16 ( .A(s44[1]), .Z(n9) );
  CMXI2X1 U17 ( .A0(n10), .A1(n9), .S(n8), .Z(sum4[3]) );
endmodule


module Add_half_6977 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6978 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3489 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6978 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6977 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6979 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6980 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3490 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6980 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6979 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6981 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6982 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3491 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6982 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6981 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6983 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6984 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3492 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6984 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6983 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_873 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3492 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3491 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3490 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3489 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out10), .A1(c_out11), .S(n4), .Z(c_out2) );
  CMXI2X1 U4 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U5 ( .A(n1), .Z(n4) );
  CIVX2 U6 ( .A(s1), .Z(n3) );
  CIVX2 U7 ( .A(s2), .Z(n2) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_6985 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6986 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3493 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6986 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6985 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6987 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6988 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3494 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6988 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6987 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6989 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_6990 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3495 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6990 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6989 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6991 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_6992 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3496 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6992 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6991 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_874 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_3496 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3495 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3494 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3493 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_6993 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6994 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3497 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6994 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6993 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6995 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6996 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3498 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6996 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6995 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6997 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_6998 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3499 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_6998 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6997 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_6999 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7000 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3500 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7000 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_6999 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_875 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8;

  Add_full_3500 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3499 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3498 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3497 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_out10), .Z(n3) );
  CIVX2 U4 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U5 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U6 ( .A(n1), .Z(n6) );
  CMXI2X1 U7 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U8 ( .A(s1), .Z(n5) );
  CIVX2 U9 ( .A(s2), .Z(n4) );
  CMXI2X1 U10 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(s3), .Z(n8) );
  CIVX2 U12 ( .A(s4), .Z(n7) );
  CMXI2X1 U13 ( .A0(n8), .A1(n7), .S(n6), .Z(sum2[1]) );
endmodule


module Add_half_7001 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7002 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3501 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7002 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7001 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7003 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7004 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3502 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7004 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7003 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7005 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7006 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3503 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7006 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7005 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7007 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7008 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3504 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7008 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7007 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_876 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3504 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3503 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3502 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3501 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_219 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_876 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_875 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_874 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_873 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2XL U3 ( .A0(s43[1]), .A1(s44[1]), .S(n4), .Z(sum4[3]) );
  CMX2XL U4 ( .A0(s43[0]), .A1(s44[0]), .S(n4), .Z(sum4[2]) );
  CMX2X1 U5 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CMX2X1 U6 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U7 ( .A(c_out410), .Z(n3) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U10 ( .A(n1), .Z(n4) );
  CMXI2X1 U11 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out4) );
endmodule


module Add_half_7009 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7010 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3505 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7010 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7009 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7011 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7012 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3506 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7012 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7011 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7013 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7014 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3507 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7014 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7013 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7015 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7016 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3508 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7016 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7015 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_877 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1;

  Add_full_3508 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3507 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3506 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3505 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_7017 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7018 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3509 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7018 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7017 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7019 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7020 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3510 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7020 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7019 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7021 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7022 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3511 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7022 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7021 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7023 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7024 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3512 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7024 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7023 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_878 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1;

  Add_full_3512 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3511 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3510 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3509 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n1), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n1), .Z(c_out2) );
  CMX2X1 U6 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_7025 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7026 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3513 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7026 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7025 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7027 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7028 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3514 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7028 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7027 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7029 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7030 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3515 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7030 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7029 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7031 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7032 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3516 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7032 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7031 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_879 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3516 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3515 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3514 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3513 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_7033 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7034 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3517 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7034 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7033 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7035 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7036 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3518 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7036 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7035 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7037 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7038 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3519 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7038 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7037 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7039 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7040 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3520 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7040 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7039 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_880 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3520 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3519 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3518 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3517 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_220 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_880 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_879 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_878 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_877 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMXI2XL U3 ( .A0(n9), .A1(n8), .S(n10), .Z(sum4[2]) );
  CIVX2 U4 ( .A(c_out410), .Z(n3) );
  CIVX2 U5 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n10) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n10), .Z(c_out4) );
  CIVX2 U9 ( .A(s41[0]), .Z(n5) );
  CIVX2 U10 ( .A(s42[0]), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U12 ( .A(s41[1]), .Z(n7) );
  CIVX2 U13 ( .A(s42[1]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U15 ( .A(s43[0]), .Z(n9) );
  CIVX2 U16 ( .A(s44[0]), .Z(n8) );
  CIVX2 U17 ( .A(s43[1]), .Z(n12) );
  CIVX2 U18 ( .A(s44[1]), .Z(n11) );
  CMXI2X1 U19 ( .A0(n12), .A1(n11), .S(n10), .Z(sum4[3]) );
endmodule


module bit8_55 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   n15, c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6,
         n7, n9, n10, n11, n12, n13, n14;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_220 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_219 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_218 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_217 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CMX2X1 U3 ( .A0(s83[3]), .A1(s84[3]), .S(n2), .Z(sum8[7]) );
  CND2X1 U4 ( .A(n6), .B(n7), .Z(sum8[0]) );
  CND2XL U5 ( .A(c_in8), .B(s82[0]), .Z(n7) );
  CNIVX4 U6 ( .A(n15), .Z(sum8[5]) );
  CNIVX1 U7 ( .A(c_in8), .Z(n1) );
  CMXI2X1 U8 ( .A0(n13), .A1(n12), .S(n2), .Z(n15) );
  CMX2X2 U9 ( .A0(s81[2]), .A1(s82[2]), .S(n1), .Z(sum8[2]) );
  CIVXL U10 ( .A(c_in8), .Z(n5) );
  CMXI2XL U11 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n3) );
  CIVXL U12 ( .A(n3), .Z(n2) );
  CMX2X2 U13 ( .A0(s81[3]), .A1(s82[3]), .S(n1), .Z(sum8[3]) );
  CIVXL U14 ( .A(n3), .Z(n4) );
  CIVX2 U15 ( .A(n9), .Z(n14) );
  CMX2XL U16 ( .A0(s81[1]), .A1(s82[1]), .S(c_in8), .Z(sum8[1]) );
  CMX2X2 U17 ( .A0(s83[2]), .A1(s84[2]), .S(n4), .Z(sum8[6]) );
  CMX2X2 U18 ( .A0(c_out810), .A1(c_out811), .S(n14), .Z(c_out8) );
  CND2X1 U19 ( .A(s81[0]), .B(n5), .Z(n6) );
  CMXI2X1 U20 ( .A0(n11), .A1(n10), .S(n14), .Z(sum8[4]) );
  CMXI2X1 U21 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n9) );
  CIVX2 U22 ( .A(s83[0]), .Z(n11) );
  CIVX2 U23 ( .A(s84[0]), .Z(n10) );
  CIVX2 U24 ( .A(s83[1]), .Z(n13) );
  CIVX2 U25 ( .A(s84[1]), .Z(n12) );
endmodule


module Add_half_7041 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7042 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3521 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7042 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7041 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7043 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7044 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3522 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7044 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7043 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7045 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_7046 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3523 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7046 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7045 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7047 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7048 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3524 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7048 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7047 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_881 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3524 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3523 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3522 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3521 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2XL U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n4) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module Add_half_7049 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7050 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3525 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7050 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7049 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7051 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7052 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3526 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7052 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7051 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7053 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_7054 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3527 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7054 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7053 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7055 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7056 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3528 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7056 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7055 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_882 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2;

  Add_full_3528 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3527 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3526 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3525 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2XL U3 ( .A0(s3), .A1(s4), .S(n2), .Z(sum2[1]) );
  CMX2XL U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CMX2X1 U5 ( .A0(c_out10), .A1(c_out11), .S(n2), .Z(c_out2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n2) );
endmodule


module Add_half_7057 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7058 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3529 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7058 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7057 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7059 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7060 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3530 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7060 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7059 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7061 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1, n2;

  CIVXL U1 ( .A(a), .Z(n1) );
  CIVXL U2 ( .A(n1), .Z(n2) );
  CEOXL U3 ( .A(b), .B(n2), .Z(sum) );
  CAN2X1 U4 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7062 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX2 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3531 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7062 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7061 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7063 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7064 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX3 U1 ( .A(b), .Z(n1) );
  CENX2 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3532 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7064 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7063 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_883 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3532 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3531 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3530 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3529 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMXI2XL U3 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
  CIVX1 U4 ( .A(n1), .Z(n4) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U10 ( .A(s3), .Z(n6) );
  CIVX2 U11 ( .A(s4), .Z(n5) );
endmodule


module Add_half_7065 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7066 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3533 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7066 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7065 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7067 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7068 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3534 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7068 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7067 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7069 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7070 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX2 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3535 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7070 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7069 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7071 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(n1), .Z(sum) );
  CNIVXL U3 ( .A(a), .Z(n1) );
endmodule


module Add_half_7072 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3536 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7072 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7071 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_884 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_3536 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3535 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3534 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3533 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U3 ( .A(c_in2), .Z(n1) );
  CIVX2 U4 ( .A(n2), .Z(n5) );
  CIVX1 U5 ( .A(c_out10), .Z(n4) );
  CMXI2X1 U6 ( .A0(c_out01), .A1(c_out00), .S(n1), .Z(n2) );
  CMX2XL U7 ( .A0(s3), .A1(s4), .S(n5), .Z(sum2[1]) );
  CMX2X1 U8 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U9 ( .A(c_out11), .Z(n3) );
  CMXI2X1 U10 ( .A0(n4), .A1(n3), .S(n5), .Z(c_out2) );
endmodule


module bit4_221 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_884 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_883 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_882 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_881 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CMX2X1 U3 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CIVXL U4 ( .A(n2), .Z(n1) );
  CMXI2X1 U5 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n2) );
  CIVX1 U6 ( .A(n2), .Z(n5) );
  CMX2XL U7 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U8 ( .A0(c_out410), .A1(c_out411), .S(n5), .Z(c_out4) );
  CMX2X1 U9 ( .A0(s41[1]), .A1(s42[1]), .S(c_in4), .Z(sum4[1]) );
  CIVX2 U10 ( .A(s41[0]), .Z(n4) );
  CIVX2 U11 ( .A(s42[0]), .Z(n3) );
  CMXI2X1 U12 ( .A0(n4), .A1(n3), .S(c_in4), .Z(sum4[0]) );
endmodule


module Add_half_7073 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7074 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3537 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7074 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7073 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7075 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7076 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3538 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7076 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7075 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7077 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7078 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3539 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7078 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7077 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7079 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7080 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3540 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7080 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7079 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module bit2_885 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3540 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3539 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3538 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3537 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CMX2X1 U3 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U4 ( .A(c_out10), .Z(n3) );
  CIVX2 U5 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U6 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U7 ( .A(n1), .Z(n4) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
  CIVX2 U9 ( .A(s3), .Z(n6) );
  CIVX2 U10 ( .A(s4), .Z(n5) );
  CMXI2X1 U11 ( .A0(n6), .A1(n5), .S(n4), .Z(sum2[1]) );
endmodule


module Add_half_7081 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U2 ( .A(b), .Z(n2) );
  CENX1 U3 ( .A(a), .B(n2), .Z(sum) );
endmodule


module Add_half_7082 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3541 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7082 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7081 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7083 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7084 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3542 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7084 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7083 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7085 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7086 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3543 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7086 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7085 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7087 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7088 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3544 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7088 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7087 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX1 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_886 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3544 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3543 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3542 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3541 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(s1), .Z(n5) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CIVX2 U8 ( .A(n1), .Z(n6) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_7089 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7090 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3545 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7090 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7089 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7091 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7092 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3546 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7092 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7091 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7093 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7094 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3547 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7094 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7093 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7095 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7096 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3548 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7096 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7095 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_887 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3548 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3547 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3546 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3545 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n6) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n6), .Z(sum2[1]) );
  CIVX2 U5 ( .A(c_out10), .Z(n3) );
  CIVX2 U6 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U7 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U8 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out2) );
  CIVX2 U9 ( .A(s1), .Z(n5) );
  CIVX2 U10 ( .A(s2), .Z(n4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_7097 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7098 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3549 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7098 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7097 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7099 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7100 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3550 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7100 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7099 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7101 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CENXL U2 ( .A(n2), .B(a), .Z(sum) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_7102 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3551 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7102 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7101 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7103 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7104 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(a), .B(b), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3552 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7104 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7103 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X1 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_888 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4;

  Add_full_3552 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3551 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3550 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3549 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX1 U3 ( .A(n1), .Z(n4) );
  CMX2XL U4 ( .A0(s3), .A1(s4), .S(n4), .Z(sum2[1]) );
  CMX2X1 U5 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U6 ( .A(c_out10), .Z(n3) );
  CIVX2 U7 ( .A(c_out11), .Z(n2) );
  CMXI2X1 U8 ( .A0(c_out00), .A1(c_out01), .S(c_in2), .Z(n1) );
  CMXI2X1 U9 ( .A0(n3), .A1(n2), .S(n4), .Z(c_out2) );
endmodule


module bit4_222 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_888 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_887 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_886 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_885 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CIVX1 U3 ( .A(c_out410), .Z(n3) );
  CIVX1 U4 ( .A(n1), .Z(n6) );
  CMX2XL U5 ( .A0(s43[1]), .A1(s44[1]), .S(n6), .Z(sum4[3]) );
  CMX2XL U6 ( .A0(s43[0]), .A1(s44[0]), .S(n6), .Z(sum4[2]) );
  CMX2X1 U7 ( .A0(s41[0]), .A1(s42[0]), .S(c_in4), .Z(sum4[0]) );
  CIVX2 U8 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U9 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n6), .Z(c_out4) );
  CIVX2 U11 ( .A(s41[1]), .Z(n5) );
  CIVX2 U12 ( .A(s42[1]), .Z(n4) );
  CMXI2X1 U13 ( .A0(n5), .A1(n4), .S(c_in4), .Z(sum4[1]) );
endmodule


module Add_half_7105 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7106 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3553 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7106 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7105 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7107 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7108 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3554 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7108 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7107 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7109 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CNIVXL U1 ( .A(a), .Z(n1) );
  CEOXL U2 ( .A(b), .B(n1), .Z(sum) );
  CAN2X1 U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7110 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3555 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7110 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7109 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7111 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_7112 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3556 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7112 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7111 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module bit2_889 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5;

  Add_full_3556 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3555 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3554 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3553 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X2 U3 ( .A(n2), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n1) );
  CMX2XL U4 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CANR2XL U5 ( .A(n2), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n3) );
  CMX2X1 U6 ( .A0(c_out11), .A1(c_out10), .S(n1), .Z(c_out2) );
  CMXI2XL U7 ( .A0(n5), .A1(n4), .S(n3), .Z(sum2[1]) );
  CIVX2 U8 ( .A(c_in2), .Z(n2) );
  CIVX2 U9 ( .A(s4), .Z(n5) );
  CIVX2 U10 ( .A(s3), .Z(n4) );
endmodule


module Add_half_7113 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_half_7114 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3557 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7114 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7113 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7115 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_7116 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3558 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7116 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7115 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7117 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7118 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(n1), .B(a), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3559 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7118 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7117 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2X2 U1 ( .A(n2), .B(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w3), .Z(n2) );
  CIVX2 U3 ( .A(w2), .Z(n1) );
endmodule


module Add_half_7119 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(a), .B(b), .Z(c_out) );
  CEOXL U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7120 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3560 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7120 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7119 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_890 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6, n7, n8, n9;

  Add_full_3560 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3559 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3558 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3557 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2X1 U3 ( .A(n3), .B(n4), .Z(c_out2) );
  CANR2X1 U4 ( .A(n6), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n1) );
  CANR2X1 U5 ( .A(n6), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n5) );
  CND2X2 U6 ( .A(c_out11), .B(n2), .Z(n3) );
  CND2X1 U7 ( .A(c_out10), .B(n5), .Z(n4) );
  CIVX2 U8 ( .A(n1), .Z(n2) );
  CIVXL U9 ( .A(s2), .Z(n7) );
  CIVX1 U10 ( .A(s1), .Z(n8) );
  CANR2XL U11 ( .A(n6), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n9) );
  CMX2XL U12 ( .A0(s4), .A1(s3), .S(n9), .Z(sum2[1]) );
  CIVX2 U13 ( .A(c_in2), .Z(n6) );
  CMXI2X1 U14 ( .A0(n8), .A1(n7), .S(c_in2), .Z(sum2[0]) );
endmodule


module Add_half_7121 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7122 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3561 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7122 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7121 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7123 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7124 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3562 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7124 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7123 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7125 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7126 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3563 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7126 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7125 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7127 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7128 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3564 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7128 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7127 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_891 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3564 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3563 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3562 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3561 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7129 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7130 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3565 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7130 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7129 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7131 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_half_7132 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3566 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7132 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7131 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7133 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7134 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3567 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7134 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7133 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7135 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7136 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3568 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7136 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7135 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_892 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3568 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3567 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3566 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3565 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_223 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_892 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_891 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_890 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_889 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n4), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n4), .Z(sum4[0]) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX1 U4 ( .A(c_out411), .Z(n2) );
  CMXI2X1 U5 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out4) );
  CIVX2 U6 ( .A(c_out410), .Z(n3) );
  CMX2X1 U7 ( .A0(s43[1]), .A1(s44[1]), .S(n1), .Z(sum4[3]) );
  CMX2X1 U10 ( .A0(s43[0]), .A1(s44[0]), .S(n1), .Z(sum4[2]) );
  CIVX2 U11 ( .A(c_in4), .Z(n4) );
endmodule


module Add_half_7137 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(n2), .B(a), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_7138 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3569 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7138 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7137 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7139 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_7140 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3570 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7140 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7139 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7141 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7142 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX2 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3571 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7142 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7141 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_7143 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7144 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3572 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7144 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7143 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module bit2_893 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3;

  Add_full_3572 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3571 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3570 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3569 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CANR2X2 U3 ( .A(n2), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n1) );
  CANR2XL U4 ( .A(n2), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n3) );
  CMX2XL U5 ( .A0(s4), .A1(s3), .S(n3), .Z(sum2[1]) );
  CMX2X1 U6 ( .A0(c_out11), .A1(c_out10), .S(n1), .Z(c_out2) );
  CMX2X1 U7 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U8 ( .A(c_in2), .Z(n2) );
endmodule


module Add_half_7145 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_7146 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3573 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7146 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7145 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7147 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n2;

  CENXL U1 ( .A(a), .B(n2), .Z(sum) );
  CAN2XL U2 ( .A(a), .B(b), .Z(c_out) );
  CIVX2 U3 ( .A(b), .Z(n2) );
endmodule


module Add_half_7148 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2XL U1 ( .A(a), .B(b), .Z(c_out) );
  CEOX1 U2 ( .A(a), .B(b), .Z(sum) );
endmodule


module Add_full_3574 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7148 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7147 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w3), .B(w2), .Z(c_out) );
endmodule


module Add_half_7149 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7150 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3575 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1, n2;

  Add_half_7150 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7149 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CIVX2 U1 ( .A(w3), .Z(n2) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
  CND2X2 U3 ( .A(n2), .B(n1), .Z(c_out) );
endmodule


module Add_half_7151 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOXL U1 ( .A(a), .B(b), .Z(sum) );
  CAN2X1 U2 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_half_7152 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;
  wire   n1;

  CIVX2 U1 ( .A(b), .Z(n1) );
  CENX1 U2 ( .A(a), .B(n1), .Z(sum) );
  CAN2XL U3 ( .A(a), .B(b), .Z(c_out) );
endmodule


module Add_full_3576 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3, n1;

  Add_half_7152 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7151 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  CND2IX1 U1 ( .B(w3), .A(n1), .Z(c_out) );
  CIVX2 U2 ( .A(w2), .Z(n1) );
endmodule


module bit2_894 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n2, n3, n4,
         n5, n6;

  Add_full_3576 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3575 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3574 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3573 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CND2X1 U3 ( .A(n2), .B(n3), .Z(c_out2) );
  CND2X2 U4 ( .A(c_out11), .B(n1), .Z(n2) );
  CND2X1 U5 ( .A(c_out10), .B(n6), .Z(n3) );
  CIVX2 U6 ( .A(n6), .Z(n1) );
  CANR2XL U7 ( .A(n5), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n4) );
  CMX2XL U8 ( .A0(s4), .A1(s3), .S(n4), .Z(sum2[1]) );
  CANR2X2 U9 ( .A(n5), .B(c_out00), .C(c_in2), .D(c_out01), .Z(n6) );
  CMX2X1 U10 ( .A0(s1), .A1(s2), .S(c_in2), .Z(sum2[0]) );
  CIVX2 U11 ( .A(c_in2), .Z(n5) );
endmodule


module Add_half_7153 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7154 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3577 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7154 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7153 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7155 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7156 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3578 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7156 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7155 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7157 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7158 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3579 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7158 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7157 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7159 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7160 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3580 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7160 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7159 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_895 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3580 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3579 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3578 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3577 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module Add_half_7161 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7162 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3581 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7162 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7161 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7163 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7164 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3582 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7164 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7163 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7165 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7166 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CAN2X1 U1 ( .A(b), .B(a), .Z(c_out) );
  CEOX1 U2 ( .A(b), .B(a), .Z(sum) );
endmodule


module Add_full_3583 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7166 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7165 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module Add_half_7167 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_half_7168 ( sum, c_out, a, b );
  input a, b;
  output sum, c_out;


  CEOX1 U1 ( .A(b), .B(a), .Z(sum) );
  CAN2X1 U2 ( .A(b), .B(a), .Z(c_out) );
endmodule


module Add_full_3584 ( sum, c_out, a, b, c_in );
  input a, b, c_in;
  output sum, c_out;
  wire   w1, w2, w3;

  Add_half_7168 M1 ( .sum(w1), .c_out(w2), .a(a), .b(b) );
  Add_half_7167 M2 ( .sum(sum), .c_out(w3), .a(w1), .b(c_in) );
  COR2X1 U1 ( .A(w2), .B(w3), .Z(c_out) );
endmodule


module bit2_896 ( sum2, c_out2, a2, b2, c_in2 );
  output [1:0] sum2;
  input [1:0] a2;
  input [1:0] b2;
  input c_in2;
  output c_out2;
  wire   s1, c_out00, s2, c_out01, s3, c_out10, s4, c_out11, n1, n4, n5;

  Add_full_3584 A1 ( .sum(s1), .c_out(c_out00), .a(a2[0]), .b(b2[0]), .c_in(
        1'b0) );
  Add_full_3583 A2 ( .sum(s2), .c_out(c_out01), .a(a2[0]), .b(b2[0]), .c_in(
        1'b1) );
  Add_full_3582 A3 ( .sum(s3), .c_out(c_out10), .a(a2[1]), .b(b2[1]), .c_in(
        1'b0) );
  Add_full_3581 A4 ( .sum(s4), .c_out(c_out11), .a(a2[1]), .b(b2[1]), .c_in(
        1'b1) );
  CIVX2 U4 ( .A(n1), .Z(n5) );
  CIVX2 U5 ( .A(c_in2), .Z(n4) );
  CAOR2X1 U6 ( .A(s4), .B(n5), .C(s3), .D(n1), .Z(sum2[1]) );
  CAOR2X1 U7 ( .A(s2), .B(c_in2), .C(s1), .D(n4), .Z(sum2[0]) );
  CAOR2X1 U8 ( .A(c_out11), .B(n5), .C(c_out10), .D(n1), .Z(c_out2) );
  CANR2X1 U3 ( .A(c_out01), .B(c_in2), .C(c_out00), .D(n4), .Z(n1) );
endmodule


module bit4_224 ( sum4, c_out4, a4, b4, c_in4 );
  output [3:0] sum4;
  input [3:0] a4;
  input [3:0] b4;
  input c_in4;
  output c_out4;
  wire   c_out400, c_out401, c_out410, c_out411, n1, n2, n3, n4, n5, n6, n7,
         n8;
  wire   [1:0] s41;
  wire   [1:0] s42;
  wire   [1:0] s43;
  wire   [1:0] s44;

  bit2_896 A41 ( .sum2(s41), .c_out2(c_out400), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b0) );
  bit2_895 A42 ( .sum2(s42), .c_out2(c_out401), .a2(a4[1:0]), .b2(b4[1:0]), 
        .c_in2(1'b1) );
  bit2_894 A43 ( .sum2(s43), .c_out2(c_out410), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b0) );
  bit2_893 A44 ( .sum2(s44), .c_out2(c_out411), .a2(a4[3:2]), .b2(b4[3:2]), 
        .c_in2(1'b1) );
  CAOR2X1 U8 ( .A(s42[1]), .B(c_in4), .C(s41[1]), .D(n8), .Z(sum4[1]) );
  CAOR2X1 U9 ( .A(s42[0]), .B(c_in4), .C(s41[0]), .D(n8), .Z(sum4[0]) );
  CMX2X1 U3 ( .A0(c_out400), .A1(c_out401), .S(c_in4), .Z(n1) );
  CIVX1 U4 ( .A(c_out411), .Z(n2) );
  CIVX2 U5 ( .A(c_out410), .Z(n3) );
  CIVX1 U6 ( .A(s44[0]), .Z(n4) );
  CIVX1 U7 ( .A(s43[0]), .Z(n5) );
  CMXI2X1 U10 ( .A0(n3), .A1(n2), .S(n1), .Z(c_out4) );
  CMXI2X1 U11 ( .A0(n5), .A1(n4), .S(n1), .Z(sum4[2]) );
  CIVX2 U12 ( .A(s43[1]), .Z(n7) );
  CIVX2 U13 ( .A(s44[1]), .Z(n6) );
  CMXI2X1 U14 ( .A0(n7), .A1(n6), .S(n1), .Z(sum4[3]) );
  CIVX2 U15 ( .A(c_in4), .Z(n8) );
endmodule


module bit8_56 ( sum8, c_out8, a8, b8, c_in8 );
  output [7:0] sum8;
  input [7:0] a8;
  input [7:0] b8;
  input c_in8;
  output c_out8;
  wire   c_out800, c_out801, c_out810, c_out811, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16;
  wire   [3:0] s81;
  wire   [3:0] s82;
  wire   [3:0] s83;
  wire   [3:0] s84;

  bit4_224 A81 ( .sum4(s81), .c_out4(c_out800), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b0) );
  bit4_223 A82 ( .sum4(s82), .c_out4(c_out801), .a4(a8[3:0]), .b4(b8[3:0]), 
        .c_in4(1'b1) );
  bit4_222 A83 ( .sum4(s83), .c_out4(c_out810), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b0) );
  bit4_221 A84 ( .sum4(s84), .c_out4(c_out811), .a4(a8[7:4]), .b4(b8[7:4]), 
        .c_in4(1'b1) );
  CAOR2X1 U12 ( .A(s82[1]), .B(c_in8), .C(s81[1]), .D(n16), .Z(sum8[1]) );
  CAOR2X1 U13 ( .A(s82[0]), .B(c_in8), .C(s81[0]), .D(n16), .Z(sum8[0]) );
  CMXI2X2 U3 ( .A0(n10), .A1(n9), .S(c_in8), .Z(sum8[3]) );
  CMXI2X1 U4 ( .A0(c_out800), .A1(c_out801), .S(c_in8), .Z(n6) );
  CIVX1 U5 ( .A(s84[2]), .Z(n11) );
  CMX2X1 U6 ( .A0(s83[0]), .A1(s84[0]), .S(n13), .Z(sum8[4]) );
  CMXI2X1 U7 ( .A0(n8), .A1(n7), .S(c_in8), .Z(sum8[2]) );
  CNIVX2 U8 ( .A(n1), .Z(n2) );
  CIVX1 U9 ( .A(s82[2]), .Z(n7) );
  CND2X1 U10 ( .A(c_out810), .B(n3), .Z(n4) );
  CND2X2 U11 ( .A(n4), .B(n5), .Z(c_out8) );
  CIVXL U14 ( .A(s84[3]), .Z(n14) );
  CIVXL U15 ( .A(n6), .Z(n1) );
  CIVX1 U16 ( .A(n6), .Z(n13) );
  CMXI2X1 U17 ( .A0(n12), .A1(n11), .S(n2), .Z(sum8[6]) );
  CIVX1 U18 ( .A(s83[3]), .Z(n15) );
  CIVX1 U19 ( .A(s83[2]), .Z(n12) );
  CND2X1 U20 ( .A(c_out811), .B(n13), .Z(n5) );
  CIVX1 U21 ( .A(n13), .Z(n3) );
  CMX2X1 U22 ( .A0(s83[1]), .A1(s84[1]), .S(n1), .Z(sum8[5]) );
  CMXI2XL U23 ( .A0(n15), .A1(n14), .S(n2), .Z(sum8[7]) );
  CIVX2 U24 ( .A(s81[2]), .Z(n8) );
  CIVX2 U25 ( .A(s81[3]), .Z(n10) );
  CIVX2 U26 ( .A(s82[3]), .Z(n9) );
  CIVX2 U27 ( .A(c_in8), .Z(n16) );
endmodule


module bit32_14 ( a32, b32, sum32, c_out32, c_in32 );
  input [31:0] a32;
  input [31:0] b32;
  output [31:0] sum32;
  input c_in32;
  output c_out32;
  wire   c1, c2, c3;

  bit8_56 A321 ( .sum8(sum32[7:0]), .c_out8(c1), .a8(a32[7:0]), .b8(b32[7:0]), 
        .c_in8(c_in32) );
  bit8_55 A322 ( .sum8(sum32[15:8]), .c_out8(c2), .a8(a32[15:8]), .b8(
        b32[15:8]), .c_in8(c1) );
  bit8_54 A323 ( .sum8(sum32[23:16]), .c_out8(c3), .a8(a32[23:16]), .b8(
        b32[23:16]), .c_in8(c2) );
  bit8_53 A324 ( .sum8(sum32[31:24]), .c_out8(c_out32), .a8(a32[31:24]), .b8(
        b32[31:24]), .c_in8(c3) );
endmodule


module array_bin ( mlier, mcand, prodt, start, reset, valid, clock );
  input [15:0] mlier;
  input [15:0] mcand;
  output [31:0] prodt;
  input start, reset, clock;
  output valid;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, net84808, net91924, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97;
  wire   [31:0] s15;
  wire   [15:0] p0;
  wire   [15:0] p1;
  wire   [15:0] p2;
  wire   [15:0] p3;
  wire   [15:0] p4;
  wire   [15:0] p5;
  wire   [15:0] p6;
  wire   [15:0] p7;
  wire   [15:0] p8;
  wire   [15:0] p9;
  wire   [15:0] p10;
  wire   [15:0] p11;
  wire   [15:0] p12;
  wire   [15:0] p13;
  wire   [15:0] p14;
  wire   [15:0] p15;
  wire   [31:0] s1;
  wire   [31:0] s2;
  wire   [31:0] s3;
  wire   [31:0] s4;
  wire   [31:0] s5;
  wire   [31:0] s6;
  wire   [31:0] s7;
  wire   [31:0] s8;
  wire   [31:0] s9;
  wire   [31:0] s10;
  wire   [31:0] s11;
  wire   [31:0] s12;
  wire   [31:0] s13;
  wire   [31:0] s14;

  bit32_0 A0 ( .a32({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, p0}), .b32({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        p1, 1'b0}), .sum32(s1), .c_in32(1'b0) );
  bit32_14 A1 ( .a32({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, p2, 1'b0, 1'b0}), .b32({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, p3, 1'b0, 
        1'b0, 1'b0}), .sum32(s2), .c_in32(1'b0) );
  bit32_13 A2 ( .a32({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, p4, 1'b0, 1'b0, 1'b0, 1'b0}), .b32({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, p5[15:3], n40, p5[1:0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum32(s3), .c_in32(1'b0) );
  bit32_12 A3 ( .a32({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, p6, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b32({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, p7, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .sum32(s4), .c_in32(1'b0) );
  bit32_11 A4 ( .a32({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, p8, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b32({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, p9, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .sum32(s5), .c_in32(1'b0) );
  bit32_10 A5 ( .a32({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, p10, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b32({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, p11, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .sum32(s6), .c_in32(1'b0) );
  bit32_9 A6 ( .a32({1'b0, 1'b0, 1'b0, 1'b0, p12, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b32({1'b0, 1'b0, 1'b0, 
        p13, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .sum32(s7), .c_in32(1'b0) );
  bit32_8 A7 ( .a32({1'b0, 1'b0, p14, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b32({1'b0, p15, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .sum32(s8), .c_in32(1'b0) );
  bit32_7 A8 ( .a32(s1), .b32({s2[31:13], n89, s2[11:8], n39, n93, s2[5:0]}), 
        .sum32(s9), .c_in32(1'b0) );
  bit32_6 A9 ( .a32(s3), .b32(s4), .sum32(s10), .c_in32(1'b0) );
  bit32_5 A10 ( .a32({s5[31:11], n83, n95, s5[8:0]}), .b32({s6[31:21], n65, 
        s6[19:17], n84, s6[15:0]}), .sum32(s11), .c_in32(1'b0) );
  bit32_4 A11 ( .a32(s7), .b32({s8[31:25], n91, s8[23:0]}), .sum32(s12), 
        .c_in32(1'b0) );
  bit32_3 A12 ( .a32({s9[31:3], n97, s9[1:0]}), .b32({s10[31:13], n42, 
        s10[11:0]}), .sum32(s13), .c_in32(1'b0) );
  bit32_2 A13 ( .a32(s11), .b32(s12), .sum32(s14), .c_in32(1'b0) );
  bit32_1 A14 ( .a32(s13), .b32(s14), .sum32(s15), .c_in32(1'b0) );
  CFD1QXL \prodt_reg[7]  ( .D(N10), .CP(clock), .Q(prodt[7]) );
  CFD1QXL \prodt_reg[6]  ( .D(N9), .CP(clock), .Q(prodt[6]) );
  CFD1QXL \prodt_reg[5]  ( .D(N8), .CP(clock), .Q(prodt[5]) );
  CFD1QXL \prodt_reg[4]  ( .D(N7), .CP(clock), .Q(prodt[4]) );
  CFD1QXL \prodt_reg[3]  ( .D(N6), .CP(clock), .Q(prodt[3]) );
  CFD1QXL \prodt_reg[2]  ( .D(N5), .CP(clock), .Q(prodt[2]) );
  CFD1QXL \prodt_reg[1]  ( .D(N4), .CP(clock), .Q(prodt[1]) );
  CFD1QXL \prodt_reg[0]  ( .D(N3), .CP(clock), .Q(prodt[0]) );
  CFD1QXL valid_reg ( .D(net84808), .CP(clock), .Q(valid) );
  CFD1QXL \prodt_reg[19]  ( .D(N22), .CP(clock), .Q(prodt[19]) );
  CFD1QXL \prodt_reg[18]  ( .D(N21), .CP(clock), .Q(prodt[18]) );
  CFD1QXL \prodt_reg[17]  ( .D(N20), .CP(clock), .Q(prodt[17]) );
  CFD1QXL \prodt_reg[16]  ( .D(N19), .CP(clock), .Q(prodt[16]) );
  CFD1QXL \prodt_reg[15]  ( .D(N18), .CP(clock), .Q(prodt[15]) );
  CFD1QXL \prodt_reg[14]  ( .D(N17), .CP(clock), .Q(prodt[14]) );
  CFD1QXL \prodt_reg[13]  ( .D(N16), .CP(clock), .Q(prodt[13]) );
  CFD1QXL \prodt_reg[12]  ( .D(N15), .CP(clock), .Q(prodt[12]) );
  CFD1QXL \prodt_reg[11]  ( .D(N14), .CP(clock), .Q(prodt[11]) );
  CFD1QXL \prodt_reg[10]  ( .D(N13), .CP(clock), .Q(prodt[10]) );
  CFD1QXL \prodt_reg[9]  ( .D(N12), .CP(clock), .Q(prodt[9]) );
  CFD1QXL \prodt_reg[8]  ( .D(N11), .CP(clock), .Q(prodt[8]) );
  CFD1QX2 \prodt_reg[30]  ( .D(N33), .CP(clock), .Q(prodt[30]) );
  CFD1QX2 \prodt_reg[26]  ( .D(N29), .CP(clock), .Q(prodt[26]) );
  CFD1QX1 \prodt_reg[27]  ( .D(N30), .CP(clock), .Q(prodt[27]) );
  CFD3QX2 \prodt_reg[31]  ( .D(N34), .CP(clock), .CD(1'b1), .SD(1'b1), .Q(
        prodt[31]) );
  CFD3QX2 \prodt_reg[29]  ( .D(N32), .CP(clock), .CD(1'b1), .SD(1'b1), .Q(
        prodt[29]) );
  CFD3QX2 \prodt_reg[28]  ( .D(N31), .CP(clock), .CD(1'b1), .SD(1'b1), .Q(
        prodt[28]) );
  CFD1QX1 \prodt_reg[25]  ( .D(N28), .CP(clock), .Q(prodt[25]) );
  CFD1QX1 \prodt_reg[23]  ( .D(N26), .CP(clock), .Q(prodt[23]) );
  CFD1QX1 \prodt_reg[22]  ( .D(N25), .CP(clock), .Q(prodt[22]) );
  CFD1QX1 \prodt_reg[21]  ( .D(N24), .CP(clock), .Q(prodt[21]) );
  CFD1QX1 \prodt_reg[20]  ( .D(N23), .CP(clock), .Q(prodt[20]) );
  CFD1QX1 \prodt_reg[24]  ( .D(N27), .CP(clock), .Q(prodt[24]) );
  CIVX4 U324 ( .A(n70), .Z(p11[1]) );
  CND2X2 U325 ( .A(mlier[3]), .B(mcand[3]), .Z(n35) );
  CIVX3 U326 ( .A(n35), .Z(p3[3]) );
  CND2X4 U327 ( .A(mlier[7]), .B(mcand[0]), .Z(n36) );
  CIVX2 U328 ( .A(n36), .Z(p7[0]) );
  CND2X4 U329 ( .A(mlier[7]), .B(mcand[2]), .Z(n37) );
  CIVX2 U330 ( .A(n37), .Z(p7[2]) );
  CND2X2 U331 ( .A(mlier[9]), .B(mcand[3]), .Z(n38) );
  CIVX3 U332 ( .A(n38), .Z(p9[3]) );
  CNIVX3 U333 ( .A(s2[7]), .Z(n39) );
  CIVX8 U334 ( .A(n45), .Z(p10[0]) );
  CIVX8 U335 ( .A(n75), .Z(p1[4]) );
  CIVX4 U336 ( .A(n81), .Z(p0[2]) );
  CIVX8 U337 ( .A(n77), .Z(p0[6]) );
  CIVX2 U338 ( .A(n73), .Z(p0[5]) );
  CIVX3 U339 ( .A(n66), .Z(p2[1]) );
  CAN2X2 U340 ( .A(mlier[0]), .B(mcand[3]), .Z(p0[3]) );
  CIVX8 U341 ( .A(n60), .Z(p5[1]) );
  CIVX3 U342 ( .A(n53), .Z(p4[2]) );
  CIVX8 U343 ( .A(n56), .Z(p9[1]) );
  CIVX4 U344 ( .A(n54), .Z(p8[2]) );
  CIVX3 U345 ( .A(n52), .Z(p8[1]) );
  CIVX3 U346 ( .A(n69), .Z(p10[2]) );
  CNR2IX1 U347 ( .B(s15[4]), .A(reset), .Z(N7) );
  CNR2IX1 U348 ( .B(s15[5]), .A(reset), .Z(N8) );
  CNR2IX1 U349 ( .B(s15[6]), .A(reset), .Z(N9) );
  CNR2IX1 U350 ( .B(s15[7]), .A(reset), .Z(N10) );
  CAN2X2 U351 ( .A(mlier[5]), .B(mcand[2]), .Z(n40) );
  CAN2X1 U352 ( .A(s15[26]), .B(net84808), .Z(N29) );
  CIVX12 U353 ( .A(mcand[0]), .Z(net91924) );
  CIVX4 U354 ( .A(s10[12]), .Z(n41) );
  CIVX8 U355 ( .A(n41), .Z(n42) );
  CAN2X2 U356 ( .A(mlier[9]), .B(mcand[5]), .Z(p9[5]) );
  CNR2X4 U357 ( .A(n43), .B(n44), .Z(p4[4]) );
  CIVX20 U358 ( .A(mlier[4]), .Z(n43) );
  CIVX20 U359 ( .A(mcand[4]), .Z(n44) );
  CND2X4 U360 ( .A(mlier[10]), .B(mcand[0]), .Z(n45) );
  CND2X4 U361 ( .A(mlier[5]), .B(mcand[3]), .Z(n46) );
  CIVX4 U362 ( .A(n46), .Z(p5[3]) );
  CND2IX1 U363 ( .B(reset), .A(s15[28]), .Z(n47) );
  CND2IX1 U364 ( .B(reset), .A(s15[29]), .Z(n48) );
  CND2IX1 U365 ( .B(reset), .A(s15[31]), .Z(n49) );
  CND2IX1 U366 ( .B(reset), .A(s15[30]), .Z(n50) );
  CIVX1 U367 ( .A(n47), .Z(N31) );
  CIVX1 U368 ( .A(n48), .Z(N32) );
  CIVX1 U369 ( .A(n49), .Z(N34) );
  CIVX1 U370 ( .A(n50), .Z(N33) );
  CIVX2 U371 ( .A(reset), .Z(net84808) );
  CND2X4 U372 ( .A(mlier[0]), .B(mcand[0]), .Z(n51) );
  CIVX8 U373 ( .A(n51), .Z(p0[0]) );
  CAN2X2 U374 ( .A(mlier[7]), .B(mcand[5]), .Z(p7[5]) );
  CAN2X2 U375 ( .A(mlier[6]), .B(mcand[6]), .Z(p6[6]) );
  CIVX2 U376 ( .A(s9[2]), .Z(n96) );
  CND2X4 U377 ( .A(mlier[9]), .B(mcand[0]), .Z(n67) );
  CAN2X2 U378 ( .A(mlier[11]), .B(mcand[3]), .Z(p11[3]) );
  CND2X4 U379 ( .A(mlier[8]), .B(mcand[1]), .Z(n52) );
  CND2X4 U380 ( .A(mlier[4]), .B(mcand[2]), .Z(n53) );
  CAN2X2 U381 ( .A(mlier[12]), .B(mcand[2]), .Z(p12[2]) );
  CAN2X2 U382 ( .A(mlier[10]), .B(mcand[1]), .Z(p10[1]) );
  CIVX8 U383 ( .A(n55), .Z(p6[2]) );
  CAN2X2 U384 ( .A(mlier[7]), .B(mcand[3]), .Z(p7[3]) );
  CAN2X2 U385 ( .A(mlier[6]), .B(mcand[4]), .Z(p6[4]) );
  CIVX8 U386 ( .A(n59), .Z(p7[1]) );
  CIVX8 U387 ( .A(n58), .Z(p4[1]) );
  CIVX8 U388 ( .A(n74), .Z(p0[1]) );
  CAN2X2 U389 ( .A(mlier[13]), .B(mcand[1]), .Z(p13[1]) );
  CAN2X2 U390 ( .A(mlier[2]), .B(mcand[6]), .Z(p2[6]) );
  CIVX8 U391 ( .A(n82), .Z(p1[1]) );
  CND2X4 U392 ( .A(mlier[8]), .B(mcand[2]), .Z(n54) );
  CAN2X2 U393 ( .A(mlier[10]), .B(mcand[3]), .Z(p10[3]) );
  CIVX8 U394 ( .A(n57), .Z(p12[0]) );
  CND2X4 U395 ( .A(mlier[5]), .B(mcand[0]), .Z(n68) );
  CND2X4 U396 ( .A(mlier[6]), .B(mcand[2]), .Z(n55) );
  CND2X4 U397 ( .A(mlier[9]), .B(mcand[1]), .Z(n56) );
  CND2X4 U398 ( .A(mlier[12]), .B(mcand[0]), .Z(n57) );
  CND2X4 U399 ( .A(mlier[4]), .B(mcand[1]), .Z(n58) );
  CND2X4 U400 ( .A(mlier[7]), .B(mcand[1]), .Z(n59) );
  CND2X4 U401 ( .A(mlier[5]), .B(mcand[1]), .Z(n60) );
  CAN2X2 U405 ( .A(mlier[6]), .B(mcand[3]), .Z(p6[3]) );
  CAN2X4 U406 ( .A(mlier[8]), .B(mcand[5]), .Z(p8[5]) );
  CAN2X4 U407 ( .A(mlier[9]), .B(mcand[4]), .Z(p9[4]) );
  CND2X4 U408 ( .A(mlier[3]), .B(mcand[0]), .Z(n72) );
  CIVX2 U409 ( .A(s6[20]), .Z(n64) );
  CIVX4 U410 ( .A(n64), .Z(n65) );
  CND2X4 U411 ( .A(mlier[2]), .B(mcand[1]), .Z(n66) );
  CAN2X2 U412 ( .A(mlier[11]), .B(mcand[2]), .Z(p11[2]) );
  CAN2X2 U413 ( .A(mlier[8]), .B(mcand[4]), .Z(p8[4]) );
  CIVX8 U414 ( .A(n72), .Z(p3[0]) );
  CIVX8 U415 ( .A(n68), .Z(p5[0]) );
  CIVX8 U416 ( .A(n67), .Z(p9[0]) );
  CAN2X2 U417 ( .A(mlier[0]), .B(mcand[8]), .Z(p0[8]) );
  CAN2X2 U418 ( .A(mlier[12]), .B(mcand[1]), .Z(p12[1]) );
  CND2X4 U419 ( .A(mlier[10]), .B(mcand[2]), .Z(n69) );
  CAN2X2 U420 ( .A(mlier[3]), .B(mcand[5]), .Z(p3[5]) );
  CND2X4 U421 ( .A(mlier[11]), .B(mcand[1]), .Z(n70) );
  CNR2X4 U422 ( .A(n71), .B(net91924), .Z(p1[0]) );
  CIVX20 U423 ( .A(mlier[1]), .Z(n71) );
  CIVX8 U424 ( .A(n78), .Z(p8[0]) );
  CND2X4 U425 ( .A(mlier[0]), .B(mcand[5]), .Z(n73) );
  CAN2X2 U426 ( .A(mlier[1]), .B(mcand[7]), .Z(p1[7]) );
  CIVX8 U427 ( .A(n86), .Z(p2[2]) );
  CND2X4 U428 ( .A(mlier[0]), .B(mcand[1]), .Z(n74) );
  CIVX8 U429 ( .A(n80), .Z(p0[4]) );
  CIVX2 U430 ( .A(s2[6]), .Z(n92) );
  CND2X4 U431 ( .A(mlier[1]), .B(mcand[4]), .Z(n75) );
  CIVX8 U432 ( .A(n76), .Z(p4[0]) );
  CIVX8 U433 ( .A(n85), .Z(p1[3]) );
  CAN2X2 U434 ( .A(mlier[6]), .B(mcand[1]), .Z(p6[1]) );
  CND2X4 U435 ( .A(mlier[4]), .B(mcand[0]), .Z(n76) );
  CIVX8 U436 ( .A(n79), .Z(p6[0]) );
  CND2X4 U437 ( .A(mlier[0]), .B(mcand[6]), .Z(n77) );
  CND2X4 U438 ( .A(mlier[8]), .B(mcand[0]), .Z(n78) );
  CAN2X2 U439 ( .A(mlier[1]), .B(mcand[5]), .Z(p1[5]) );
  CND2X4 U440 ( .A(mlier[6]), .B(mcand[0]), .Z(n79) );
  CND2X4 U441 ( .A(mlier[0]), .B(mcand[4]), .Z(n80) );
  CND2X4 U442 ( .A(mlier[0]), .B(mcand[2]), .Z(n81) );
  CND2X4 U443 ( .A(mlier[1]), .B(mcand[1]), .Z(n82) );
  CNIVX4 U444 ( .A(s5[10]), .Z(n83) );
  CNIVX4 U445 ( .A(s6[16]), .Z(n84) );
  CAN2X2 U446 ( .A(mlier[11]), .B(mcand[0]), .Z(p11[0]) );
  CAN2X2 U447 ( .A(mlier[13]), .B(mcand[0]), .Z(p13[0]) );
  CND2X4 U448 ( .A(mlier[1]), .B(mcand[3]), .Z(n85) );
  CAN2X2 U449 ( .A(mlier[2]), .B(mcand[4]), .Z(p2[4]) );
  CAN2X4 U450 ( .A(mlier[2]), .B(mcand[3]), .Z(p2[3]) );
  CAN2X4 U451 ( .A(mlier[3]), .B(mcand[2]), .Z(p3[2]) );
  CIVX8 U452 ( .A(n88), .Z(p2[0]) );
  CIVX8 U453 ( .A(n87), .Z(p3[1]) );
  CND2X4 U454 ( .A(mlier[2]), .B(mcand[2]), .Z(n86) );
  CND2X4 U455 ( .A(mlier[3]), .B(mcand[1]), .Z(n87) );
  CND2X4 U456 ( .A(mlier[2]), .B(mcand[0]), .Z(n88) );
  CAN2X2 U457 ( .A(mlier[15]), .B(mcand[0]), .Z(p15[0]) );
  CAN2X2 U458 ( .A(mcand[0]), .B(mlier[14]), .Z(p14[0]) );
  CAN2X2 U459 ( .A(mlier[1]), .B(mcand[2]), .Z(p1[2]) );
  CNIVX4 U460 ( .A(s2[12]), .Z(n89) );
  CAN2X1 U461 ( .A(mlier[3]), .B(mcand[4]), .Z(p3[4]) );
  CAN2X1 U462 ( .A(mlier[4]), .B(mcand[3]), .Z(p4[3]) );
  CAN2X1 U463 ( .A(mlier[2]), .B(mcand[5]), .Z(p2[5]) );
  CAN2X1 U464 ( .A(mlier[9]), .B(mcand[2]), .Z(p9[2]) );
  CAN2X1 U465 ( .A(mlier[8]), .B(mcand[3]), .Z(p8[3]) );
  CAN2X1 U466 ( .A(mlier[13]), .B(mcand[2]), .Z(p13[2]) );
  CAN2X1 U467 ( .A(mcand[1]), .B(mlier[14]), .Z(p14[1]) );
  CAN2X1 U468 ( .A(mlier[12]), .B(mcand[3]), .Z(p12[3]) );
  CAN2X1 U469 ( .A(mcand[2]), .B(mlier[14]), .Z(p14[2]) );
  CAN2X1 U470 ( .A(mlier[15]), .B(mcand[1]), .Z(p15[1]) );
  CIVX4 U471 ( .A(n92), .Z(n93) );
  CIVX4 U472 ( .A(n94), .Z(n95) );
  CIVX4 U473 ( .A(n90), .Z(n91) );
  CAN2X1 U474 ( .A(mcand[3]), .B(mlier[14]), .Z(p14[3]) );
  CAN2X1 U475 ( .A(mlier[8]), .B(mcand[7]), .Z(p8[7]) );
  CAN2X1 U476 ( .A(mlier[15]), .B(mcand[2]), .Z(p15[2]) );
  CAN2X1 U477 ( .A(mlier[9]), .B(mcand[6]), .Z(p9[6]) );
  CAN2X1 U478 ( .A(mlier[10]), .B(mcand[4]), .Z(p10[4]) );
  CAN2X1 U479 ( .A(mcand[4]), .B(mlier[14]), .Z(p14[4]) );
  CIVX4 U480 ( .A(n96), .Z(n97) );
  CAN2X1 U481 ( .A(mlier[12]), .B(mcand[5]), .Z(p12[5]) );
  CAN2X1 U482 ( .A(mlier[13]), .B(mcand[4]), .Z(p13[4]) );
  CNR2IX1 U483 ( .B(s15[1]), .A(reset), .Z(N4) );
  CNR2IX1 U484 ( .B(s15[2]), .A(reset), .Z(N5) );
  CNR2IX1 U485 ( .B(s15[3]), .A(reset), .Z(N6) );
  CNR2IX1 U486 ( .B(s15[0]), .A(reset), .Z(N3) );
  CIVX2 U487 ( .A(s8[24]), .Z(n90) );
  CIVX2 U488 ( .A(s5[9]), .Z(n94) );
  CAN2X1 U489 ( .A(s15[8]), .B(net84808), .Z(N11) );
  CAN2X1 U490 ( .A(s15[9]), .B(net84808), .Z(N12) );
  CAN2X1 U491 ( .A(s15[10]), .B(net84808), .Z(N13) );
  CAN2X1 U492 ( .A(s15[11]), .B(net84808), .Z(N14) );
  CAN2X1 U493 ( .A(s15[12]), .B(net84808), .Z(N15) );
  CAN2X1 U494 ( .A(s15[13]), .B(net84808), .Z(N16) );
  CAN2X1 U495 ( .A(s15[14]), .B(net84808), .Z(N17) );
  CAN2X1 U496 ( .A(s15[15]), .B(net84808), .Z(N18) );
  CAN2X1 U497 ( .A(s15[16]), .B(net84808), .Z(N19) );
  CAN2X1 U498 ( .A(s15[17]), .B(net84808), .Z(N20) );
  CAN2X1 U499 ( .A(s15[18]), .B(net84808), .Z(N21) );
  CAN2X1 U500 ( .A(s15[19]), .B(net84808), .Z(N22) );
  CAN2X1 U501 ( .A(s15[20]), .B(net84808), .Z(N23) );
  CAN2X1 U502 ( .A(s15[21]), .B(net84808), .Z(N24) );
  CAN2X1 U503 ( .A(s15[22]), .B(net84808), .Z(N25) );
  CAN2X1 U504 ( .A(s15[23]), .B(net84808), .Z(N26) );
  CAN2X1 U505 ( .A(s15[24]), .B(net84808), .Z(N27) );
  CAN2X1 U506 ( .A(s15[25]), .B(net84808), .Z(N28) );
  CAN2X1 U507 ( .A(s15[27]), .B(net84808), .Z(N30) );
  CAN2X1 U508 ( .A(mlier[14]), .B(mcand[15]), .Z(p14[15]) );
  CAN2X1 U509 ( .A(mcand[14]), .B(mlier[14]), .Z(p14[14]) );
  CAN2X1 U510 ( .A(mcand[13]), .B(mlier[14]), .Z(p14[13]) );
  CAN2X1 U511 ( .A(mcand[12]), .B(mlier[14]), .Z(p14[12]) );
  CAN2X1 U512 ( .A(mcand[11]), .B(mlier[14]), .Z(p14[11]) );
  CAN2X1 U513 ( .A(mcand[10]), .B(mlier[14]), .Z(p14[10]) );
  CAN2X1 U514 ( .A(mcand[9]), .B(mlier[14]), .Z(p14[9]) );
  CAN2X1 U515 ( .A(mcand[8]), .B(mlier[14]), .Z(p14[8]) );
  CAN2X1 U516 ( .A(mcand[7]), .B(mlier[14]), .Z(p14[7]) );
  CAN2X1 U517 ( .A(mcand[6]), .B(mlier[14]), .Z(p14[6]) );
  CAN2X1 U518 ( .A(mcand[5]), .B(mlier[14]), .Z(p14[5]) );
  CAN2X1 U519 ( .A(mlier[15]), .B(mcand[15]), .Z(p15[15]) );
  CAN2X1 U520 ( .A(mlier[15]), .B(mcand[14]), .Z(p15[14]) );
  CAN2X1 U521 ( .A(mlier[15]), .B(mcand[13]), .Z(p15[13]) );
  CAN2X1 U522 ( .A(mlier[15]), .B(mcand[12]), .Z(p15[12]) );
  CAN2X1 U523 ( .A(mlier[15]), .B(mcand[11]), .Z(p15[11]) );
  CAN2X1 U524 ( .A(mlier[15]), .B(mcand[10]), .Z(p15[10]) );
  CAN2X1 U525 ( .A(mlier[15]), .B(mcand[9]), .Z(p15[9]) );
  CAN2X1 U526 ( .A(mlier[15]), .B(mcand[8]), .Z(p15[8]) );
  CAN2X1 U527 ( .A(mlier[15]), .B(mcand[7]), .Z(p15[7]) );
  CAN2X1 U528 ( .A(mlier[15]), .B(mcand[6]), .Z(p15[6]) );
  CAN2X1 U529 ( .A(mlier[15]), .B(mcand[5]), .Z(p15[5]) );
  CAN2X1 U530 ( .A(mlier[15]), .B(mcand[4]), .Z(p15[4]) );
  CAN2X1 U531 ( .A(mlier[15]), .B(mcand[3]), .Z(p15[3]) );
  CAN2X1 U532 ( .A(mlier[12]), .B(mcand[15]), .Z(p12[15]) );
  CAN2X1 U533 ( .A(mlier[12]), .B(mcand[14]), .Z(p12[14]) );
  CAN2X1 U534 ( .A(mlier[12]), .B(mcand[13]), .Z(p12[13]) );
  CAN2X1 U535 ( .A(mlier[12]), .B(mcand[12]), .Z(p12[12]) );
  CAN2X1 U536 ( .A(mlier[12]), .B(mcand[11]), .Z(p12[11]) );
  CAN2X1 U537 ( .A(mlier[12]), .B(mcand[10]), .Z(p12[10]) );
  CAN2X1 U538 ( .A(mlier[12]), .B(mcand[9]), .Z(p12[9]) );
  CAN2X1 U539 ( .A(mlier[12]), .B(mcand[8]), .Z(p12[8]) );
  CAN2X1 U540 ( .A(mlier[12]), .B(mcand[7]), .Z(p12[7]) );
  CAN2X1 U541 ( .A(mlier[12]), .B(mcand[6]), .Z(p12[6]) );
  CAN2X1 U542 ( .A(mlier[12]), .B(mcand[4]), .Z(p12[4]) );
  CAN2X1 U543 ( .A(mlier[13]), .B(mcand[15]), .Z(p13[15]) );
  CAN2X1 U544 ( .A(mlier[13]), .B(mcand[14]), .Z(p13[14]) );
  CAN2X1 U545 ( .A(mlier[13]), .B(mcand[13]), .Z(p13[13]) );
  CAN2X1 U546 ( .A(mlier[13]), .B(mcand[12]), .Z(p13[12]) );
  CAN2X1 U547 ( .A(mlier[13]), .B(mcand[11]), .Z(p13[11]) );
  CAN2X1 U548 ( .A(mlier[13]), .B(mcand[10]), .Z(p13[10]) );
  CAN2X1 U549 ( .A(mlier[13]), .B(mcand[9]), .Z(p13[9]) );
  CAN2X1 U550 ( .A(mlier[13]), .B(mcand[8]), .Z(p13[8]) );
  CAN2X1 U551 ( .A(mlier[13]), .B(mcand[7]), .Z(p13[7]) );
  CAN2X1 U552 ( .A(mlier[13]), .B(mcand[6]), .Z(p13[6]) );
  CAN2X1 U553 ( .A(mlier[13]), .B(mcand[5]), .Z(p13[5]) );
  CAN2X1 U554 ( .A(mlier[13]), .B(mcand[3]), .Z(p13[3]) );
  CAN2X1 U555 ( .A(mlier[10]), .B(mcand[15]), .Z(p10[15]) );
  CAN2X1 U556 ( .A(mlier[10]), .B(mcand[14]), .Z(p10[14]) );
  CAN2X1 U557 ( .A(mlier[10]), .B(mcand[13]), .Z(p10[13]) );
  CAN2X1 U558 ( .A(mlier[10]), .B(mcand[12]), .Z(p10[12]) );
  CAN2X1 U559 ( .A(mlier[10]), .B(mcand[11]), .Z(p10[11]) );
  CAN2X1 U560 ( .A(mlier[10]), .B(mcand[10]), .Z(p10[10]) );
  CAN2X1 U561 ( .A(mlier[10]), .B(mcand[9]), .Z(p10[9]) );
  CAN2X1 U562 ( .A(mlier[10]), .B(mcand[8]), .Z(p10[8]) );
  CAN2X1 U563 ( .A(mlier[10]), .B(mcand[7]), .Z(p10[7]) );
  CAN2X1 U564 ( .A(mlier[10]), .B(mcand[6]), .Z(p10[6]) );
  CAN2X1 U565 ( .A(mlier[10]), .B(mcand[5]), .Z(p10[5]) );
  CAN2X1 U566 ( .A(mlier[11]), .B(mcand[15]), .Z(p11[15]) );
  CAN2X1 U567 ( .A(mlier[11]), .B(mcand[14]), .Z(p11[14]) );
  CAN2X1 U568 ( .A(mlier[11]), .B(mcand[13]), .Z(p11[13]) );
  CAN2X1 U569 ( .A(mlier[11]), .B(mcand[12]), .Z(p11[12]) );
  CAN2X1 U570 ( .A(mlier[11]), .B(mcand[11]), .Z(p11[11]) );
  CAN2X1 U571 ( .A(mlier[11]), .B(mcand[10]), .Z(p11[10]) );
  CAN2X1 U572 ( .A(mlier[11]), .B(mcand[9]), .Z(p11[9]) );
  CAN2X1 U573 ( .A(mlier[11]), .B(mcand[8]), .Z(p11[8]) );
  CAN2X1 U574 ( .A(mlier[11]), .B(mcand[7]), .Z(p11[7]) );
  CAN2X1 U575 ( .A(mlier[11]), .B(mcand[6]), .Z(p11[6]) );
  CAN2X1 U576 ( .A(mlier[11]), .B(mcand[5]), .Z(p11[5]) );
  CAN2X1 U577 ( .A(mlier[11]), .B(mcand[4]), .Z(p11[4]) );
  CAN2X1 U578 ( .A(mlier[8]), .B(mcand[15]), .Z(p8[15]) );
  CAN2X1 U579 ( .A(mlier[8]), .B(mcand[14]), .Z(p8[14]) );
  CAN2X1 U580 ( .A(mlier[8]), .B(mcand[13]), .Z(p8[13]) );
  CAN2X1 U581 ( .A(mlier[8]), .B(mcand[12]), .Z(p8[12]) );
  CAN2X1 U582 ( .A(mlier[8]), .B(mcand[11]), .Z(p8[11]) );
  CAN2X1 U583 ( .A(mlier[8]), .B(mcand[10]), .Z(p8[10]) );
  CAN2X1 U584 ( .A(mlier[8]), .B(mcand[9]), .Z(p8[9]) );
  CAN2X1 U585 ( .A(mlier[8]), .B(mcand[8]), .Z(p8[8]) );
  CAN2X1 U586 ( .A(mlier[8]), .B(mcand[6]), .Z(p8[6]) );
  CAN2X1 U587 ( .A(mlier[9]), .B(mcand[15]), .Z(p9[15]) );
  CAN2X1 U588 ( .A(mlier[9]), .B(mcand[14]), .Z(p9[14]) );
  CAN2X1 U589 ( .A(mlier[9]), .B(mcand[13]), .Z(p9[13]) );
  CAN2X1 U590 ( .A(mlier[9]), .B(mcand[12]), .Z(p9[12]) );
  CAN2X1 U591 ( .A(mlier[9]), .B(mcand[11]), .Z(p9[11]) );
  CAN2X1 U592 ( .A(mlier[9]), .B(mcand[10]), .Z(p9[10]) );
  CAN2X1 U593 ( .A(mlier[9]), .B(mcand[9]), .Z(p9[9]) );
  CAN2X1 U594 ( .A(mlier[9]), .B(mcand[8]), .Z(p9[8]) );
  CAN2X1 U595 ( .A(mlier[9]), .B(mcand[7]), .Z(p9[7]) );
  CAN2X1 U596 ( .A(mlier[6]), .B(mcand[15]), .Z(p6[15]) );
  CAN2X1 U597 ( .A(mlier[6]), .B(mcand[14]), .Z(p6[14]) );
  CAN2X1 U598 ( .A(mlier[6]), .B(mcand[13]), .Z(p6[13]) );
  CAN2X1 U599 ( .A(mlier[6]), .B(mcand[12]), .Z(p6[12]) );
  CAN2X1 U600 ( .A(mlier[6]), .B(mcand[11]), .Z(p6[11]) );
  CAN2X1 U601 ( .A(mlier[6]), .B(mcand[10]), .Z(p6[10]) );
  CAN2X1 U602 ( .A(mlier[6]), .B(mcand[9]), .Z(p6[9]) );
  CAN2X1 U603 ( .A(mlier[6]), .B(mcand[8]), .Z(p6[8]) );
  CAN2X1 U604 ( .A(mlier[6]), .B(mcand[7]), .Z(p6[7]) );
  CAN2X1 U605 ( .A(mlier[6]), .B(mcand[5]), .Z(p6[5]) );
  CAN2X1 U606 ( .A(mlier[7]), .B(mcand[15]), .Z(p7[15]) );
  CAN2X1 U607 ( .A(mlier[7]), .B(mcand[14]), .Z(p7[14]) );
  CAN2X1 U608 ( .A(mlier[7]), .B(mcand[13]), .Z(p7[13]) );
  CAN2X1 U609 ( .A(mlier[7]), .B(mcand[12]), .Z(p7[12]) );
  CAN2X1 U610 ( .A(mlier[7]), .B(mcand[11]), .Z(p7[11]) );
  CAN2X1 U611 ( .A(mlier[7]), .B(mcand[10]), .Z(p7[10]) );
  CAN2X1 U612 ( .A(mlier[7]), .B(mcand[9]), .Z(p7[9]) );
  CAN2X1 U613 ( .A(mlier[7]), .B(mcand[8]), .Z(p7[8]) );
  CAN2X1 U614 ( .A(mlier[7]), .B(mcand[7]), .Z(p7[7]) );
  CAN2X1 U615 ( .A(mlier[7]), .B(mcand[6]), .Z(p7[6]) );
  CAN2X1 U616 ( .A(mlier[7]), .B(mcand[4]), .Z(p7[4]) );
  CAN2X1 U617 ( .A(mlier[4]), .B(mcand[15]), .Z(p4[15]) );
  CAN2X1 U618 ( .A(mlier[4]), .B(mcand[14]), .Z(p4[14]) );
  CAN2X1 U619 ( .A(mlier[4]), .B(mcand[13]), .Z(p4[13]) );
  CAN2X1 U620 ( .A(mlier[4]), .B(mcand[12]), .Z(p4[12]) );
  CAN2X1 U621 ( .A(mlier[4]), .B(mcand[11]), .Z(p4[11]) );
  CAN2X1 U622 ( .A(mlier[4]), .B(mcand[10]), .Z(p4[10]) );
  CAN2X1 U623 ( .A(mlier[4]), .B(mcand[9]), .Z(p4[9]) );
  CAN2X1 U624 ( .A(mlier[4]), .B(mcand[8]), .Z(p4[8]) );
  CAN2X1 U625 ( .A(mlier[4]), .B(mcand[7]), .Z(p4[7]) );
  CAN2X1 U626 ( .A(mlier[4]), .B(mcand[6]), .Z(p4[6]) );
  CAN2X1 U627 ( .A(mlier[4]), .B(mcand[5]), .Z(p4[5]) );
  CAN2X1 U628 ( .A(mlier[5]), .B(mcand[15]), .Z(p5[15]) );
  CAN2X1 U629 ( .A(mlier[5]), .B(mcand[14]), .Z(p5[14]) );
  CAN2X1 U630 ( .A(mlier[5]), .B(mcand[13]), .Z(p5[13]) );
  CAN2X1 U631 ( .A(mlier[5]), .B(mcand[12]), .Z(p5[12]) );
  CAN2X1 U632 ( .A(mlier[5]), .B(mcand[11]), .Z(p5[11]) );
  CAN2X1 U633 ( .A(mlier[5]), .B(mcand[10]), .Z(p5[10]) );
  CAN2X1 U634 ( .A(mlier[5]), .B(mcand[9]), .Z(p5[9]) );
  CAN2X1 U635 ( .A(mlier[5]), .B(mcand[8]), .Z(p5[8]) );
  CAN2X1 U636 ( .A(mlier[5]), .B(mcand[7]), .Z(p5[7]) );
  CAN2X1 U637 ( .A(mlier[5]), .B(mcand[6]), .Z(p5[6]) );
  CAN2X1 U638 ( .A(mlier[5]), .B(mcand[5]), .Z(p5[5]) );
  CAN2X1 U639 ( .A(mlier[5]), .B(mcand[4]), .Z(p5[4]) );
  CAN2X1 U640 ( .A(mlier[2]), .B(mcand[15]), .Z(p2[15]) );
  CAN2X1 U641 ( .A(mlier[2]), .B(mcand[14]), .Z(p2[14]) );
  CAN2X1 U642 ( .A(mlier[2]), .B(mcand[13]), .Z(p2[13]) );
  CAN2X1 U643 ( .A(mlier[2]), .B(mcand[12]), .Z(p2[12]) );
  CAN2X1 U644 ( .A(mlier[2]), .B(mcand[11]), .Z(p2[11]) );
  CAN2X1 U645 ( .A(mlier[2]), .B(mcand[10]), .Z(p2[10]) );
  CAN2X1 U646 ( .A(mlier[2]), .B(mcand[9]), .Z(p2[9]) );
  CAN2X1 U647 ( .A(mlier[2]), .B(mcand[8]), .Z(p2[8]) );
  CAN2X1 U648 ( .A(mlier[2]), .B(mcand[7]), .Z(p2[7]) );
  CAN2X1 U649 ( .A(mlier[3]), .B(mcand[15]), .Z(p3[15]) );
  CAN2X1 U650 ( .A(mlier[3]), .B(mcand[14]), .Z(p3[14]) );
  CAN2X1 U651 ( .A(mlier[3]), .B(mcand[13]), .Z(p3[13]) );
  CAN2X1 U652 ( .A(mlier[3]), .B(mcand[12]), .Z(p3[12]) );
  CAN2X1 U653 ( .A(mlier[3]), .B(mcand[11]), .Z(p3[11]) );
  CAN2X1 U654 ( .A(mlier[3]), .B(mcand[10]), .Z(p3[10]) );
  CAN2X1 U655 ( .A(mlier[3]), .B(mcand[9]), .Z(p3[9]) );
  CAN2X1 U656 ( .A(mlier[3]), .B(mcand[8]), .Z(p3[8]) );
  CAN2X1 U657 ( .A(mlier[3]), .B(mcand[7]), .Z(p3[7]) );
  CAN2X1 U658 ( .A(mlier[3]), .B(mcand[6]), .Z(p3[6]) );
  CAN2X1 U659 ( .A(mlier[0]), .B(mcand[15]), .Z(p0[15]) );
  CAN2X1 U660 ( .A(mlier[0]), .B(mcand[14]), .Z(p0[14]) );
  CAN2X1 U661 ( .A(mlier[0]), .B(mcand[13]), .Z(p0[13]) );
  CAN2X1 U662 ( .A(mlier[0]), .B(mcand[12]), .Z(p0[12]) );
  CAN2X1 U663 ( .A(mlier[0]), .B(mcand[11]), .Z(p0[11]) );
  CAN2X1 U664 ( .A(mlier[0]), .B(mcand[10]), .Z(p0[10]) );
  CAN2X1 U665 ( .A(mlier[0]), .B(mcand[9]), .Z(p0[9]) );
  CAN2X1 U666 ( .A(mlier[0]), .B(mcand[7]), .Z(p0[7]) );
  CAN2X1 U667 ( .A(mlier[1]), .B(mcand[15]), .Z(p1[15]) );
  CAN2X1 U668 ( .A(mlier[1]), .B(mcand[14]), .Z(p1[14]) );
  CAN2X1 U669 ( .A(mlier[1]), .B(mcand[13]), .Z(p1[13]) );
  CAN2X1 U670 ( .A(mlier[1]), .B(mcand[12]), .Z(p1[12]) );
  CAN2X1 U671 ( .A(mlier[1]), .B(mcand[11]), .Z(p1[11]) );
  CAN2X1 U672 ( .A(mlier[1]), .B(mcand[10]), .Z(p1[10]) );
  CAN2X1 U673 ( .A(mlier[1]), .B(mcand[9]), .Z(p1[9]) );
  CAN2X1 U674 ( .A(mlier[1]), .B(mcand[8]), .Z(p1[8]) );
  CAN2X1 U675 ( .A(mlier[1]), .B(mcand[6]), .Z(p1[6]) );
endmodule

